// Developed by: Amir Yazdanbakhsh
// Email: a.yazdanbakhsh@gatech.edu

`timescale 1ns/1ps
module asin_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000000000000000010000; // input=0.00048828125, output=0.000488281269403
			11'd1: out = 32'b00000000000000000000000000110000; // input=0.00146484375, output=0.00146484427387
			11'd2: out = 32'b00000000000000000000000001010000; // input=0.00244140625, output=0.00244140867533
			11'd3: out = 32'b00000000000000000000000001110000; // input=0.00341796875, output=0.00341797540511
			11'd4: out = 32'b00000000000000000000000010010000; // input=0.00439453125, output=0.00439454539458
			11'd5: out = 32'b00000000000000000000000010110000; // input=0.00537109375, output=0.00537111957513
			11'd6: out = 32'b00000000000000000000000011010000; // input=0.00634765625, output=0.00634769887818
			11'd7: out = 32'b00000000000000000000000011110000; // input=0.00732421875, output=0.0073242842352
			11'd8: out = 32'b00000000000000000000000100010000; // input=0.00830078125, output=0.0083008765777
			11'd9: out = 32'b00000000000000000000000100110000; // input=0.00927734375, output=0.00927747683727
			11'd10: out = 32'b00000000000000000000000101010000; // input=0.01025390625, output=0.0102540859456
			11'd11: out = 32'b00000000000000000000000101110000; // input=0.01123046875, output=0.0112307048343
			11'd12: out = 32'b00000000000000000000000110010000; // input=0.01220703125, output=0.0122073344352
			11'd13: out = 32'b00000000000000000000000110110000; // input=0.01318359375, output=0.0131839756803
			11'd14: out = 32'b00000000000000000000000111010000; // input=0.01416015625, output=0.0141606295016
			11'd15: out = 32'b00000000000000000000000111110000; // input=0.01513671875, output=0.0151372968311
			11'd16: out = 32'b00000000000000000000001000010000; // input=0.01611328125, output=0.016113978601
			11'd17: out = 32'b00000000000000000000001000110000; // input=0.01708984375, output=0.0170906757438
			11'd18: out = 32'b00000000000000000000001001010000; // input=0.01806640625, output=0.0180673891919
			11'd19: out = 32'b00000000000000000000001001110000; // input=0.01904296875, output=0.0190441198779
			11'd20: out = 32'b00000000000000000000001010010000; // input=0.02001953125, output=0.0200208687346
			11'd21: out = 32'b00000000000000000000001010110000; // input=0.02099609375, output=0.0209976366949
			11'd22: out = 32'b00000000000000000000001011010000; // input=0.02197265625, output=0.0219744246919
			11'd23: out = 32'b00000000000000000000001011110000; // input=0.02294921875, output=0.0229512336589
			11'd24: out = 32'b00000000000000000000001100010000; // input=0.02392578125, output=0.0239280645293
			11'd25: out = 32'b00000000000000000000001100110000; // input=0.02490234375, output=0.0249049182366
			11'd26: out = 32'b00000000000000000000001101010000; // input=0.02587890625, output=0.0258817957149
			11'd27: out = 32'b00000000000000000000001101110000; // input=0.02685546875, output=0.026858697898
			11'd28: out = 32'b00000000000000000000001110010000; // input=0.02783203125, output=0.0278356257202
			11'd29: out = 32'b00000000000000000000001110110000; // input=0.02880859375, output=0.028812580116
			11'd30: out = 32'b00000000000000000000001111010000; // input=0.02978515625, output=0.0297895620201
			11'd31: out = 32'b00000000000000000000001111110000; // input=0.03076171875, output=0.0307665723674
			11'd32: out = 32'b00000000000000000000010000010000; // input=0.03173828125, output=0.0317436120931
			11'd33: out = 32'b00000000000000000000010000110000; // input=0.03271484375, output=0.0327206821325
			11'd34: out = 32'b00000000000000000000010001010000; // input=0.03369140625, output=0.0336977834215
			11'd35: out = 32'b00000000000000000000010001110000; // input=0.03466796875, output=0.0346749168959
			11'd36: out = 32'b00000000000000000000010010010000; // input=0.03564453125, output=0.0356520834919
			11'd37: out = 32'b00000000000000000000010010110000; // input=0.03662109375, output=0.0366292841462
			11'd38: out = 32'b00000000000000000000010011010000; // input=0.03759765625, output=0.0376065197954
			11'd39: out = 32'b00000000000000000000010011110000; // input=0.03857421875, output=0.0385837913767
			11'd40: out = 32'b00000000000000000000010100010000; // input=0.03955078125, output=0.0395610998276
			11'd41: out = 32'b00000000000000000000010100110000; // input=0.04052734375, output=0.0405384460857
			11'd42: out = 32'b00000000000000000000010101010000; // input=0.04150390625, output=0.0415158310892
			11'd43: out = 32'b00000000000000000000010101110000; // input=0.04248046875, output=0.0424932557764
			11'd44: out = 32'b00000000000000000000010110010000; // input=0.04345703125, output=0.0434707210861
			11'd45: out = 32'b00000000000000000000010110110000; // input=0.04443359375, output=0.0444482279573
			11'd46: out = 32'b00000000000000000000010111010001; // input=0.04541015625, output=0.0454257773296
			11'd47: out = 32'b00000000000000000000010111110001; // input=0.04638671875, output=0.0464033701426
			11'd48: out = 32'b00000000000000000000011000010001; // input=0.04736328125, output=0.0473810073367
			11'd49: out = 32'b00000000000000000000011000110001; // input=0.04833984375, output=0.0483586898524
			11'd50: out = 32'b00000000000000000000011001010001; // input=0.04931640625, output=0.0493364186307
			11'd51: out = 32'b00000000000000000000011001110001; // input=0.05029296875, output=0.0503141946129
			11'd52: out = 32'b00000000000000000000011010010001; // input=0.05126953125, output=0.0512920187407
			11'd53: out = 32'b00000000000000000000011010110001; // input=0.05224609375, output=0.0522698919565
			11'd54: out = 32'b00000000000000000000011011010001; // input=0.05322265625, output=0.0532478152028
			11'd55: out = 32'b00000000000000000000011011110001; // input=0.05419921875, output=0.0542257894226
			11'd56: out = 32'b00000000000000000000011100010001; // input=0.05517578125, output=0.0552038155595
			11'd57: out = 32'b00000000000000000000011100110001; // input=0.05615234375, output=0.0561818945573
			11'd58: out = 32'b00000000000000000000011101010001; // input=0.05712890625, output=0.0571600273605
			11'd59: out = 32'b00000000000000000000011101110001; // input=0.05810546875, output=0.0581382149139
			11'd60: out = 32'b00000000000000000000011110010001; // input=0.05908203125, output=0.0591164581629
			11'd61: out = 32'b00000000000000000000011110110001; // input=0.06005859375, output=0.0600947580532
			11'd62: out = 32'b00000000000000000000011111010001; // input=0.06103515625, output=0.0610731155313
			11'd63: out = 32'b00000000000000000000011111110001; // input=0.06201171875, output=0.0620515315438
			11'd64: out = 32'b00000000000000000000100000010001; // input=0.06298828125, output=0.0630300070381
			11'd65: out = 32'b00000000000000000000100000110001; // input=0.06396484375, output=0.064008542962
			11'd66: out = 32'b00000000000000000000100001010001; // input=0.06494140625, output=0.064987140264
			11'd67: out = 32'b00000000000000000000100001110010; // input=0.06591796875, output=0.0659657998927
			11'd68: out = 32'b00000000000000000000100010010010; // input=0.06689453125, output=0.0669445227978
			11'd69: out = 32'b00000000000000000000100010110010; // input=0.06787109375, output=0.0679233099292
			11'd70: out = 32'b00000000000000000000100011010010; // input=0.06884765625, output=0.0689021622373
			11'd71: out = 32'b00000000000000000000100011110010; // input=0.06982421875, output=0.0698810806733
			11'd72: out = 32'b00000000000000000000100100010010; // input=0.07080078125, output=0.070860066189
			11'd73: out = 32'b00000000000000000000100100110010; // input=0.07177734375, output=0.0718391197364
			11'd74: out = 32'b00000000000000000000100101010010; // input=0.07275390625, output=0.0728182422686
			11'd75: out = 32'b00000000000000000000100101110010; // input=0.07373046875, output=0.0737974347388
			11'd76: out = 32'b00000000000000000000100110010010; // input=0.07470703125, output=0.0747766981013
			11'd77: out = 32'b00000000000000000000100110110010; // input=0.07568359375, output=0.0757560333106
			11'd78: out = 32'b00000000000000000000100111010010; // input=0.07666015625, output=0.0767354413221
			11'd79: out = 32'b00000000000000000000100111110011; // input=0.07763671875, output=0.0777149230917
			11'd80: out = 32'b00000000000000000000101000010011; // input=0.07861328125, output=0.0786944795761
			11'd81: out = 32'b00000000000000000000101000110011; // input=0.07958984375, output=0.0796741117323
			11'd82: out = 32'b00000000000000000000101001010011; // input=0.08056640625, output=0.0806538205183
			11'd83: out = 32'b00000000000000000000101001110011; // input=0.08154296875, output=0.0816336068927
			11'd84: out = 32'b00000000000000000000101010010011; // input=0.08251953125, output=0.0826134718148
			11'd85: out = 32'b00000000000000000000101010110011; // input=0.08349609375, output=0.0835934162443
			11'd86: out = 32'b00000000000000000000101011010011; // input=0.08447265625, output=0.084573441142
			11'd87: out = 32'b00000000000000000000101011110011; // input=0.08544921875, output=0.0855535474692
			11'd88: out = 32'b00000000000000000000101100010100; // input=0.08642578125, output=0.086533736188
			11'd89: out = 32'b00000000000000000000101100110100; // input=0.08740234375, output=0.087514008261
			11'd90: out = 32'b00000000000000000000101101010100; // input=0.08837890625, output=0.0884943646517
			11'd91: out = 32'b00000000000000000000101101110100; // input=0.08935546875, output=0.0894748063244
			11'd92: out = 32'b00000000000000000000101110010100; // input=0.09033203125, output=0.0904553342441
			11'd93: out = 32'b00000000000000000000101110110100; // input=0.09130859375, output=0.0914359493765
			11'd94: out = 32'b00000000000000000000101111010100; // input=0.09228515625, output=0.0924166526881
			11'd95: out = 32'b00000000000000000000101111110100; // input=0.09326171875, output=0.0933974451461
			11'd96: out = 32'b00000000000000000000110000010101; // input=0.09423828125, output=0.0943783277186
			11'd97: out = 32'b00000000000000000000110000110101; // input=0.09521484375, output=0.0953593013745
			11'd98: out = 32'b00000000000000000000110001010101; // input=0.09619140625, output=0.0963403670833
			11'd99: out = 32'b00000000000000000000110001110101; // input=0.09716796875, output=0.0973215258156
			11'd100: out = 32'b00000000000000000000110010010101; // input=0.09814453125, output=0.0983027785426
			11'd101: out = 32'b00000000000000000000110010110101; // input=0.09912109375, output=0.0992841262364
			11'd102: out = 32'b00000000000000000000110011010110; // input=0.10009765625, output=0.10026556987
			11'd103: out = 32'b00000000000000000000110011110110; // input=0.10107421875, output=0.101247110417
			11'd104: out = 32'b00000000000000000000110100010110; // input=0.10205078125, output=0.102228748852
			11'd105: out = 32'b00000000000000000000110100110110; // input=0.10302734375, output=0.103210486151
			11'd106: out = 32'b00000000000000000000110101010110; // input=0.10400390625, output=0.10419232329
			11'd107: out = 32'b00000000000000000000110101110110; // input=0.10498046875, output=0.105174261246
			11'd108: out = 32'b00000000000000000000110110010111; // input=0.10595703125, output=0.106156300998
			11'd109: out = 32'b00000000000000000000110110110111; // input=0.10693359375, output=0.107138443524
			11'd110: out = 32'b00000000000000000000110111010111; // input=0.10791015625, output=0.108120689804
			11'd111: out = 32'b00000000000000000000110111110111; // input=0.10888671875, output=0.10910304082
			11'd112: out = 32'b00000000000000000000111000010111; // input=0.10986328125, output=0.110085497553
			11'd113: out = 32'b00000000000000000000111000110111; // input=0.11083984375, output=0.111068060986
			11'd114: out = 32'b00000000000000000000111001011000; // input=0.11181640625, output=0.112050732102
			11'd115: out = 32'b00000000000000000000111001111000; // input=0.11279296875, output=0.113033511886
			11'd116: out = 32'b00000000000000000000111010011000; // input=0.11376953125, output=0.114016401324
			11'd117: out = 32'b00000000000000000000111010111000; // input=0.11474609375, output=0.114999401402
			11'd118: out = 32'b00000000000000000000111011011001; // input=0.11572265625, output=0.115982513109
			11'd119: out = 32'b00000000000000000000111011111001; // input=0.11669921875, output=0.116965737431
			11'd120: out = 32'b00000000000000000000111100011001; // input=0.11767578125, output=0.11794907536
			11'd121: out = 32'b00000000000000000000111100111001; // input=0.11865234375, output=0.118932527885
			11'd122: out = 32'b00000000000000000000111101011001; // input=0.11962890625, output=0.119916095998
			11'd123: out = 32'b00000000000000000000111101111010; // input=0.12060546875, output=0.120899780692
			11'd124: out = 32'b00000000000000000000111110011010; // input=0.12158203125, output=0.12188358296
			11'd125: out = 32'b00000000000000000000111110111010; // input=0.12255859375, output=0.122867503798
			11'd126: out = 32'b00000000000000000000111111011010; // input=0.12353515625, output=0.1238515442
			11'd127: out = 32'b00000000000000000000111111111011; // input=0.12451171875, output=0.124835705164
			11'd128: out = 32'b00000000000000000001000000011011; // input=0.12548828125, output=0.125819987687
			11'd129: out = 32'b00000000000000000001000000111011; // input=0.12646484375, output=0.126804392769
			11'd130: out = 32'b00000000000000000001000001011011; // input=0.12744140625, output=0.12778892141
			11'd131: out = 32'b00000000000000000001000001111100; // input=0.12841796875, output=0.12877357461
			11'd132: out = 32'b00000000000000000001000010011100; // input=0.12939453125, output=0.129758353373
			11'd133: out = 32'b00000000000000000001000010111100; // input=0.13037109375, output=0.130743258701
			11'd134: out = 32'b00000000000000000001000011011100; // input=0.13134765625, output=0.1317282916
			11'd135: out = 32'b00000000000000000001000011111101; // input=0.13232421875, output=0.132713453074
			11'd136: out = 32'b00000000000000000001000100011101; // input=0.13330078125, output=0.133698744131
			11'd137: out = 32'b00000000000000000001000100111101; // input=0.13427734375, output=0.134684165779
			11'd138: out = 32'b00000000000000000001000101011110; // input=0.13525390625, output=0.135669719027
			11'd139: out = 32'b00000000000000000001000101111110; // input=0.13623046875, output=0.136655404886
			11'd140: out = 32'b00000000000000000001000110011110; // input=0.13720703125, output=0.137641224367
			11'd141: out = 32'b00000000000000000001000110111111; // input=0.13818359375, output=0.138627178482
			11'd142: out = 32'b00000000000000000001000111011111; // input=0.13916015625, output=0.139613268246
			11'd143: out = 32'b00000000000000000001000111111111; // input=0.14013671875, output=0.140599494675
			11'd144: out = 32'b00000000000000000001001000011111; // input=0.14111328125, output=0.141585858784
			11'd145: out = 32'b00000000000000000001001001000000; // input=0.14208984375, output=0.142572361592
			11'd146: out = 32'b00000000000000000001001001100000; // input=0.14306640625, output=0.143559004117
			11'd147: out = 32'b00000000000000000001001010000000; // input=0.14404296875, output=0.144545787379
			11'd148: out = 32'b00000000000000000001001010100001; // input=0.14501953125, output=0.145532712401
			11'd149: out = 32'b00000000000000000001001011000001; // input=0.14599609375, output=0.146519780204
			11'd150: out = 32'b00000000000000000001001011100010; // input=0.14697265625, output=0.147506991814
			11'd151: out = 32'b00000000000000000001001100000010; // input=0.14794921875, output=0.148494348255
			11'd152: out = 32'b00000000000000000001001100100010; // input=0.14892578125, output=0.149481850554
			11'd153: out = 32'b00000000000000000001001101000011; // input=0.14990234375, output=0.15046949974
			11'd154: out = 32'b00000000000000000001001101100011; // input=0.15087890625, output=0.151457296841
			11'd155: out = 32'b00000000000000000001001110000011; // input=0.15185546875, output=0.152445242889
			11'd156: out = 32'b00000000000000000001001110100100; // input=0.15283203125, output=0.153433338915
			11'd157: out = 32'b00000000000000000001001111000100; // input=0.15380859375, output=0.154421585953
			11'd158: out = 32'b00000000000000000001001111100100; // input=0.15478515625, output=0.155409985038
			11'd159: out = 32'b00000000000000000001010000000101; // input=0.15576171875, output=0.156398537206
			11'd160: out = 32'b00000000000000000001010000100101; // input=0.15673828125, output=0.157387243495
			11'd161: out = 32'b00000000000000000001010001000110; // input=0.15771484375, output=0.158376104944
			11'd162: out = 32'b00000000000000000001010001100110; // input=0.15869140625, output=0.159365122593
			11'd163: out = 32'b00000000000000000001010010000110; // input=0.15966796875, output=0.160354297484
			11'd164: out = 32'b00000000000000000001010010100111; // input=0.16064453125, output=0.161343630661
			11'd165: out = 32'b00000000000000000001010011000111; // input=0.16162109375, output=0.162333123168
			11'd166: out = 32'b00000000000000000001010011101000; // input=0.16259765625, output=0.163322776052
			11'd167: out = 32'b00000000000000000001010100001000; // input=0.16357421875, output=0.16431259036
			11'd168: out = 32'b00000000000000000001010100101001; // input=0.16455078125, output=0.165302567142
			11'd169: out = 32'b00000000000000000001010101001001; // input=0.16552734375, output=0.166292707448
			11'd170: out = 32'b00000000000000000001010101101010; // input=0.16650390625, output=0.167283012331
			11'd171: out = 32'b00000000000000000001010110001010; // input=0.16748046875, output=0.168273482845
			11'd172: out = 32'b00000000000000000001010110101010; // input=0.16845703125, output=0.169264120044
			11'd173: out = 32'b00000000000000000001010111001011; // input=0.16943359375, output=0.170254924986
			11'd174: out = 32'b00000000000000000001010111101011; // input=0.17041015625, output=0.171245898729
			11'd175: out = 32'b00000000000000000001011000001100; // input=0.17138671875, output=0.172237042333
			11'd176: out = 32'b00000000000000000001011000101100; // input=0.17236328125, output=0.173228356859
			11'd177: out = 32'b00000000000000000001011001001101; // input=0.17333984375, output=0.174219843372
			11'd178: out = 32'b00000000000000000001011001101101; // input=0.17431640625, output=0.175211502934
			11'd179: out = 32'b00000000000000000001011010001110; // input=0.17529296875, output=0.176203336613
			11'd180: out = 32'b00000000000000000001011010101110; // input=0.17626953125, output=0.177195345477
			11'd181: out = 32'b00000000000000000001011011001111; // input=0.17724609375, output=0.178187530595
			11'd182: out = 32'b00000000000000000001011011101111; // input=0.17822265625, output=0.179179893039
			11'd183: out = 32'b00000000000000000001011100010000; // input=0.17919921875, output=0.180172433881
			11'd184: out = 32'b00000000000000000001011100110000; // input=0.18017578125, output=0.181165154197
			11'd185: out = 32'b00000000000000000001011101010001; // input=0.18115234375, output=0.182158055061
			11'd186: out = 32'b00000000000000000001011101110001; // input=0.18212890625, output=0.183151137553
			11'd187: out = 32'b00000000000000000001011110010010; // input=0.18310546875, output=0.184144402751
			11'd188: out = 32'b00000000000000000001011110110011; // input=0.18408203125, output=0.185137851738
			11'd189: out = 32'b00000000000000000001011111010011; // input=0.18505859375, output=0.186131485596
			11'd190: out = 32'b00000000000000000001011111110100; // input=0.18603515625, output=0.187125305409
			11'd191: out = 32'b00000000000000000001100000010100; // input=0.18701171875, output=0.188119312266
			11'd192: out = 32'b00000000000000000001100000110101; // input=0.18798828125, output=0.189113507254
			11'd193: out = 32'b00000000000000000001100001010101; // input=0.18896484375, output=0.190107891462
			11'd194: out = 32'b00000000000000000001100001110110; // input=0.18994140625, output=0.191102465984
			11'd195: out = 32'b00000000000000000001100010010111; // input=0.19091796875, output=0.192097231912
			11'd196: out = 32'b00000000000000000001100010110111; // input=0.19189453125, output=0.193092190343
			11'd197: out = 32'b00000000000000000001100011011000; // input=0.19287109375, output=0.194087342373
			11'd198: out = 32'b00000000000000000001100011111000; // input=0.19384765625, output=0.195082689101
			11'd199: out = 32'b00000000000000000001100100011001; // input=0.19482421875, output=0.19607823163
			11'd200: out = 32'b00000000000000000001100100111010; // input=0.19580078125, output=0.19707397106
			11'd201: out = 32'b00000000000000000001100101011010; // input=0.19677734375, output=0.198069908498
			11'd202: out = 32'b00000000000000000001100101111011; // input=0.19775390625, output=0.19906604505
			11'd203: out = 32'b00000000000000000001100110011100; // input=0.19873046875, output=0.200062381825
			11'd204: out = 32'b00000000000000000001100110111100; // input=0.19970703125, output=0.201058919932
			11'd205: out = 32'b00000000000000000001100111011101; // input=0.20068359375, output=0.202055660484
			11'd206: out = 32'b00000000000000000001100111111110; // input=0.20166015625, output=0.203052604596
			11'd207: out = 32'b00000000000000000001101000011110; // input=0.20263671875, output=0.204049753384
			11'd208: out = 32'b00000000000000000001101000111111; // input=0.20361328125, output=0.205047107966
			11'd209: out = 32'b00000000000000000001101001100000; // input=0.20458984375, output=0.206044669461
			11'd210: out = 32'b00000000000000000001101010000000; // input=0.20556640625, output=0.207042438993
			11'd211: out = 32'b00000000000000000001101010100001; // input=0.20654296875, output=0.208040417685
			11'd212: out = 32'b00000000000000000001101011000010; // input=0.20751953125, output=0.209038606664
			11'd213: out = 32'b00000000000000000001101011100010; // input=0.20849609375, output=0.210037007058
			11'd214: out = 32'b00000000000000000001101100000011; // input=0.20947265625, output=0.211035619996
			11'd215: out = 32'b00000000000000000001101100100100; // input=0.21044921875, output=0.212034446612
			11'd216: out = 32'b00000000000000000001101101000101; // input=0.21142578125, output=0.21303348804
			11'd217: out = 32'b00000000000000000001101101100101; // input=0.21240234375, output=0.214032745416
			11'd218: out = 32'b00000000000000000001101110000110; // input=0.21337890625, output=0.215032219878
			11'd219: out = 32'b00000000000000000001101110100111; // input=0.21435546875, output=0.216031912567
			11'd220: out = 32'b00000000000000000001101111001000; // input=0.21533203125, output=0.217031824626
			11'd221: out = 32'b00000000000000000001101111101000; // input=0.21630859375, output=0.218031957201
			11'd222: out = 32'b00000000000000000001110000001001; // input=0.21728515625, output=0.219032311437
			11'd223: out = 32'b00000000000000000001110000101010; // input=0.21826171875, output=0.220032888484
			11'd224: out = 32'b00000000000000000001110001001011; // input=0.21923828125, output=0.221033689493
			11'd225: out = 32'b00000000000000000001110001101100; // input=0.22021484375, output=0.222034715618
			11'd226: out = 32'b00000000000000000001110010001100; // input=0.22119140625, output=0.223035968015
			11'd227: out = 32'b00000000000000000001110010101101; // input=0.22216796875, output=0.224037447841
			11'd228: out = 32'b00000000000000000001110011001110; // input=0.22314453125, output=0.225039156258
			11'd229: out = 32'b00000000000000000001110011101111; // input=0.22412109375, output=0.226041094426
			11'd230: out = 32'b00000000000000000001110100010000; // input=0.22509765625, output=0.227043263512
			11'd231: out = 32'b00000000000000000001110100110001; // input=0.22607421875, output=0.228045664681
			11'd232: out = 32'b00000000000000000001110101010001; // input=0.22705078125, output=0.229048299103
			11'd233: out = 32'b00000000000000000001110101110010; // input=0.22802734375, output=0.23005116795
			11'd234: out = 32'b00000000000000000001110110010011; // input=0.22900390625, output=0.231054272395
			11'd235: out = 32'b00000000000000000001110110110100; // input=0.22998046875, output=0.232057613615
			11'd236: out = 32'b00000000000000000001110111010101; // input=0.23095703125, output=0.233061192788
			11'd237: out = 32'b00000000000000000001110111110110; // input=0.23193359375, output=0.234065011095
			11'd238: out = 32'b00000000000000000001111000010111; // input=0.23291015625, output=0.23506906972
			11'd239: out = 32'b00000000000000000001111000111000; // input=0.23388671875, output=0.236073369847
			11'd240: out = 32'b00000000000000000001111001011001; // input=0.23486328125, output=0.237077912665
			11'd241: out = 32'b00000000000000000001111001111001; // input=0.23583984375, output=0.238082699365
			11'd242: out = 32'b00000000000000000001111010011010; // input=0.23681640625, output=0.239087731139
			11'd243: out = 32'b00000000000000000001111010111011; // input=0.23779296875, output=0.240093009183
			11'd244: out = 32'b00000000000000000001111011011100; // input=0.23876953125, output=0.241098534694
			11'd245: out = 32'b00000000000000000001111011111101; // input=0.23974609375, output=0.242104308872
			11'd246: out = 32'b00000000000000000001111100011110; // input=0.24072265625, output=0.243110332922
			11'd247: out = 32'b00000000000000000001111100111111; // input=0.24169921875, output=0.244116608046
			11'd248: out = 32'b00000000000000000001111101100000; // input=0.24267578125, output=0.245123135455
			11'd249: out = 32'b00000000000000000001111110000001; // input=0.24365234375, output=0.246129916357
			11'd250: out = 32'b00000000000000000001111110100010; // input=0.24462890625, output=0.247136951966
			11'd251: out = 32'b00000000000000000001111111000011; // input=0.24560546875, output=0.248144243497
			11'd252: out = 32'b00000000000000000001111111100100; // input=0.24658203125, output=0.249151792168
			11'd253: out = 32'b00000000000000000010000000000101; // input=0.24755859375, output=0.2501595992
			11'd254: out = 32'b00000000000000000010000000100110; // input=0.24853515625, output=0.251167665816
			11'd255: out = 32'b00000000000000000010000001000111; // input=0.24951171875, output=0.252175993242
			11'd256: out = 32'b00000000000000000010000001101000; // input=0.25048828125, output=0.253184582706
			11'd257: out = 32'b00000000000000000010000010001001; // input=0.25146484375, output=0.25419343544
			11'd258: out = 32'b00000000000000000010000010101010; // input=0.25244140625, output=0.255202552678
			11'd259: out = 32'b00000000000000000010000011001100; // input=0.25341796875, output=0.256211935655
			11'd260: out = 32'b00000000000000000010000011101101; // input=0.25439453125, output=0.257221585612
			11'd261: out = 32'b00000000000000000010000100001110; // input=0.25537109375, output=0.25823150379
			11'd262: out = 32'b00000000000000000010000100101111; // input=0.25634765625, output=0.259241691435
			11'd263: out = 32'b00000000000000000010000101010000; // input=0.25732421875, output=0.260252149793
			11'd264: out = 32'b00000000000000000010000101110001; // input=0.25830078125, output=0.261262880115
			11'd265: out = 32'b00000000000000000010000110010010; // input=0.25927734375, output=0.262273883654
			11'd266: out = 32'b00000000000000000010000110110011; // input=0.26025390625, output=0.263285161666
			11'd267: out = 32'b00000000000000000010000111010100; // input=0.26123046875, output=0.26429671541
			11'd268: out = 32'b00000000000000000010000111110110; // input=0.26220703125, output=0.265308546147
			11'd269: out = 32'b00000000000000000010001000010111; // input=0.26318359375, output=0.266320655141
			11'd270: out = 32'b00000000000000000010001000111000; // input=0.26416015625, output=0.267333043661
			11'd271: out = 32'b00000000000000000010001001011001; // input=0.26513671875, output=0.268345712975
			11'd272: out = 32'b00000000000000000010001001111010; // input=0.26611328125, output=0.269358664358
			11'd273: out = 32'b00000000000000000010001010011100; // input=0.26708984375, output=0.270371899086
			11'd274: out = 32'b00000000000000000010001010111101; // input=0.26806640625, output=0.271385418436
			11'd275: out = 32'b00000000000000000010001011011110; // input=0.26904296875, output=0.272399223693
			11'd276: out = 32'b00000000000000000010001011111111; // input=0.27001953125, output=0.273413316139
			11'd277: out = 32'b00000000000000000010001100100000; // input=0.27099609375, output=0.274427697064
			11'd278: out = 32'b00000000000000000010001101000010; // input=0.27197265625, output=0.275442367758
			11'd279: out = 32'b00000000000000000010001101100011; // input=0.27294921875, output=0.276457329516
			11'd280: out = 32'b00000000000000000010001110000100; // input=0.27392578125, output=0.277472583634
			11'd281: out = 32'b00000000000000000010001110100101; // input=0.27490234375, output=0.278488131412
			11'd282: out = 32'b00000000000000000010001111000111; // input=0.27587890625, output=0.279503974155
			11'd283: out = 32'b00000000000000000010001111101000; // input=0.27685546875, output=0.280520113167
			11'd284: out = 32'b00000000000000000010010000001001; // input=0.27783203125, output=0.28153654976
			11'd285: out = 32'b00000000000000000010010000101011; // input=0.27880859375, output=0.282553285244
			11'd286: out = 32'b00000000000000000010010001001100; // input=0.27978515625, output=0.283570320937
			11'd287: out = 32'b00000000000000000010010001101101; // input=0.28076171875, output=0.284587658157
			11'd288: out = 32'b00000000000000000010010010001111; // input=0.28173828125, output=0.285605298226
			11'd289: out = 32'b00000000000000000010010010110000; // input=0.28271484375, output=0.28662324247
			11'd290: out = 32'b00000000000000000010010011010001; // input=0.28369140625, output=0.287641492218
			11'd291: out = 32'b00000000000000000010010011110011; // input=0.28466796875, output=0.288660048801
			11'd292: out = 32'b00000000000000000010010100010100; // input=0.28564453125, output=0.289678913555
			11'd293: out = 32'b00000000000000000010010100110110; // input=0.28662109375, output=0.290698087817
			11'd294: out = 32'b00000000000000000010010101010111; // input=0.28759765625, output=0.291717572931
			11'd295: out = 32'b00000000000000000010010101111000; // input=0.28857421875, output=0.292737370241
			11'd296: out = 32'b00000000000000000010010110011010; // input=0.28955078125, output=0.293757481095
			11'd297: out = 32'b00000000000000000010010110111011; // input=0.29052734375, output=0.294777906847
			11'd298: out = 32'b00000000000000000010010111011101; // input=0.29150390625, output=0.29579864885
			11'd299: out = 32'b00000000000000000010010111111110; // input=0.29248046875, output=0.296819708463
			11'd300: out = 32'b00000000000000000010011000100000; // input=0.29345703125, output=0.29784108705
			11'd301: out = 32'b00000000000000000010011001000001; // input=0.29443359375, output=0.298862785975
			11'd302: out = 32'b00000000000000000010011001100011; // input=0.29541015625, output=0.299884806608
			11'd303: out = 32'b00000000000000000010011010000100; // input=0.29638671875, output=0.300907150321
			11'd304: out = 32'b00000000000000000010011010100110; // input=0.29736328125, output=0.30192981849
			11'd305: out = 32'b00000000000000000010011011000111; // input=0.29833984375, output=0.302952812495
			11'd306: out = 32'b00000000000000000010011011101001; // input=0.29931640625, output=0.30397613372
			11'd307: out = 32'b00000000000000000010011100001010; // input=0.30029296875, output=0.304999783551
			11'd308: out = 32'b00000000000000000010011100101100; // input=0.30126953125, output=0.306023763378
			11'd309: out = 32'b00000000000000000010011101001101; // input=0.30224609375, output=0.307048074597
			11'd310: out = 32'b00000000000000000010011101101111; // input=0.30322265625, output=0.308072718603
			11'd311: out = 32'b00000000000000000010011110010001; // input=0.30419921875, output=0.309097696799
			11'd312: out = 32'b00000000000000000010011110110010; // input=0.30517578125, output=0.310123010591
			11'd313: out = 32'b00000000000000000010011111010100; // input=0.30615234375, output=0.311148661385
			11'd314: out = 32'b00000000000000000010011111110101; // input=0.30712890625, output=0.312174650596
			11'd315: out = 32'b00000000000000000010100000010111; // input=0.30810546875, output=0.31320097964
			11'd316: out = 32'b00000000000000000010100000111001; // input=0.30908203125, output=0.314227649936
			11'd317: out = 32'b00000000000000000010100001011010; // input=0.31005859375, output=0.315254662909
			11'd318: out = 32'b00000000000000000010100001111100; // input=0.31103515625, output=0.316282019985
			11'd319: out = 32'b00000000000000000010100010011110; // input=0.31201171875, output=0.317309722597
			11'd320: out = 32'b00000000000000000010100010111111; // input=0.31298828125, output=0.318337772181
			11'd321: out = 32'b00000000000000000010100011100001; // input=0.31396484375, output=0.319366170175
			11'd322: out = 32'b00000000000000000010100100000011; // input=0.31494140625, output=0.320394918022
			11'd323: out = 32'b00000000000000000010100100100100; // input=0.31591796875, output=0.32142401717
			11'd324: out = 32'b00000000000000000010100101000110; // input=0.31689453125, output=0.32245346907
			11'd325: out = 32'b00000000000000000010100101101000; // input=0.31787109375, output=0.323483275177
			11'd326: out = 32'b00000000000000000010100110001010; // input=0.31884765625, output=0.32451343695
			11'd327: out = 32'b00000000000000000010100110101011; // input=0.31982421875, output=0.325543955852
			11'd328: out = 32'b00000000000000000010100111001101; // input=0.32080078125, output=0.326574833351
			11'd329: out = 32'b00000000000000000010100111101111; // input=0.32177734375, output=0.327606070917
			11'd330: out = 32'b00000000000000000010101000010001; // input=0.32275390625, output=0.328637670026
			11'd331: out = 32'b00000000000000000010101000110011; // input=0.32373046875, output=0.329669632158
			11'd332: out = 32'b00000000000000000010101001010100; // input=0.32470703125, output=0.330701958797
			11'd333: out = 32'b00000000000000000010101001110110; // input=0.32568359375, output=0.331734651429
			11'd334: out = 32'b00000000000000000010101010011000; // input=0.32666015625, output=0.332767711548
			11'd335: out = 32'b00000000000000000010101010111010; // input=0.32763671875, output=0.333801140649
			11'd336: out = 32'b00000000000000000010101011011100; // input=0.32861328125, output=0.334834940233
			11'd337: out = 32'b00000000000000000010101011111110; // input=0.32958984375, output=0.335869111804
			11'd338: out = 32'b00000000000000000010101100100000; // input=0.33056640625, output=0.336903656873
			11'd339: out = 32'b00000000000000000010101101000010; // input=0.33154296875, output=0.337938576951
			11'd340: out = 32'b00000000000000000010101101100011; // input=0.33251953125, output=0.338973873558
			11'd341: out = 32'b00000000000000000010101110000101; // input=0.33349609375, output=0.340009548215
			11'd342: out = 32'b00000000000000000010101110100111; // input=0.33447265625, output=0.341045602449
			11'd343: out = 32'b00000000000000000010101111001001; // input=0.33544921875, output=0.34208203779
			11'd344: out = 32'b00000000000000000010101111101011; // input=0.33642578125, output=0.343118855775
			11'd345: out = 32'b00000000000000000010110000001101; // input=0.33740234375, output=0.344156057942
			11'd346: out = 32'b00000000000000000010110000101111; // input=0.33837890625, output=0.345193645838
			11'd347: out = 32'b00000000000000000010110001010001; // input=0.33935546875, output=0.346231621009
			11'd348: out = 32'b00000000000000000010110001110011; // input=0.34033203125, output=0.347269985011
			11'd349: out = 32'b00000000000000000010110010010101; // input=0.34130859375, output=0.348308739401
			11'd350: out = 32'b00000000000000000010110010110111; // input=0.34228515625, output=0.349347885742
			11'd351: out = 32'b00000000000000000010110011011001; // input=0.34326171875, output=0.350387425601
			11'd352: out = 32'b00000000000000000010110011111100; // input=0.34423828125, output=0.351427360551
			11'd353: out = 32'b00000000000000000010110100011110; // input=0.34521484375, output=0.352467692167
			11'd354: out = 32'b00000000000000000010110101000000; // input=0.34619140625, output=0.353508422032
			11'd355: out = 32'b00000000000000000010110101100010; // input=0.34716796875, output=0.354549551733
			11'd356: out = 32'b00000000000000000010110110000100; // input=0.34814453125, output=0.355591082858
			11'd357: out = 32'b00000000000000000010110110100110; // input=0.34912109375, output=0.356633017006
			11'd358: out = 32'b00000000000000000010110111001000; // input=0.35009765625, output=0.357675355776
			11'd359: out = 32'b00000000000000000010110111101010; // input=0.35107421875, output=0.358718100774
			11'd360: out = 32'b00000000000000000010111000001101; // input=0.35205078125, output=0.359761253611
			11'd361: out = 32'b00000000000000000010111000101111; // input=0.35302734375, output=0.360804815901
			11'd362: out = 32'b00000000000000000010111001010001; // input=0.35400390625, output=0.361848789265
			11'd363: out = 32'b00000000000000000010111001110011; // input=0.35498046875, output=0.362893175329
			11'd364: out = 32'b00000000000000000010111010010110; // input=0.35595703125, output=0.363937975722
			11'd365: out = 32'b00000000000000000010111010111000; // input=0.35693359375, output=0.364983192081
			11'd366: out = 32'b00000000000000000010111011011010; // input=0.35791015625, output=0.366028826045
			11'd367: out = 32'b00000000000000000010111011111100; // input=0.35888671875, output=0.367074879261
			11'd368: out = 32'b00000000000000000010111100011111; // input=0.35986328125, output=0.368121353378
			11'd369: out = 32'b00000000000000000010111101000001; // input=0.36083984375, output=0.369168250053
			11'd370: out = 32'b00000000000000000010111101100011; // input=0.36181640625, output=0.370215570947
			11'd371: out = 32'b00000000000000000010111110000110; // input=0.36279296875, output=0.371263317726
			11'd372: out = 32'b00000000000000000010111110101000; // input=0.36376953125, output=0.372311492062
			11'd373: out = 32'b00000000000000000010111111001010; // input=0.36474609375, output=0.373360095631
			11'd374: out = 32'b00000000000000000010111111101101; // input=0.36572265625, output=0.374409130116
			11'd375: out = 32'b00000000000000000011000000001111; // input=0.36669921875, output=0.375458597205
			11'd376: out = 32'b00000000000000000011000000110001; // input=0.36767578125, output=0.37650849859
			11'd377: out = 32'b00000000000000000011000001010100; // input=0.36865234375, output=0.377558835969
			11'd378: out = 32'b00000000000000000011000001110110; // input=0.36962890625, output=0.378609611047
			11'd379: out = 32'b00000000000000000011000010011001; // input=0.37060546875, output=0.379660825532
			11'd380: out = 32'b00000000000000000011000010111011; // input=0.37158203125, output=0.38071248114
			11'd381: out = 32'b00000000000000000011000011011110; // input=0.37255859375, output=0.381764579591
			11'd382: out = 32'b00000000000000000011000100000000; // input=0.37353515625, output=0.38281712261
			11'd383: out = 32'b00000000000000000011000100100011; // input=0.37451171875, output=0.38387011193
			11'd384: out = 32'b00000000000000000011000101000101; // input=0.37548828125, output=0.384923549288
			11'd385: out = 32'b00000000000000000011000101101000; // input=0.37646484375, output=0.385977436426
			11'd386: out = 32'b00000000000000000011000110001010; // input=0.37744140625, output=0.387031775094
			11'd387: out = 32'b00000000000000000011000110101101; // input=0.37841796875, output=0.388086567045
			11'd388: out = 32'b00000000000000000011000111001111; // input=0.37939453125, output=0.38914181404
			11'd389: out = 32'b00000000000000000011000111110010; // input=0.38037109375, output=0.390197517845
			11'd390: out = 32'b00000000000000000011001000010101; // input=0.38134765625, output=0.391253680232
			11'd391: out = 32'b00000000000000000011001000110111; // input=0.38232421875, output=0.392310302978
			11'd392: out = 32'b00000000000000000011001001011010; // input=0.38330078125, output=0.393367387867
			11'd393: out = 32'b00000000000000000011001001111101; // input=0.38427734375, output=0.394424936689
			11'd394: out = 32'b00000000000000000011001010011111; // input=0.38525390625, output=0.395482951241
			11'd395: out = 32'b00000000000000000011001011000010; // input=0.38623046875, output=0.396541433322
			11'd396: out = 32'b00000000000000000011001011100101; // input=0.38720703125, output=0.397600384742
			11'd397: out = 32'b00000000000000000011001100000111; // input=0.38818359375, output=0.398659807314
			11'd398: out = 32'b00000000000000000011001100101010; // input=0.38916015625, output=0.399719702858
			11'd399: out = 32'b00000000000000000011001101001101; // input=0.39013671875, output=0.400780073201
			11'd400: out = 32'b00000000000000000011001101110000; // input=0.39111328125, output=0.401840920174
			11'd401: out = 32'b00000000000000000011001110010010; // input=0.39208984375, output=0.402902245618
			11'd402: out = 32'b00000000000000000011001110110101; // input=0.39306640625, output=0.403964051377
			11'd403: out = 32'b00000000000000000011001111011000; // input=0.39404296875, output=0.405026339302
			11'd404: out = 32'b00000000000000000011001111111011; // input=0.39501953125, output=0.406089111252
			11'd405: out = 32'b00000000000000000011010000011110; // input=0.39599609375, output=0.40715236909
			11'd406: out = 32'b00000000000000000011010001000000; // input=0.39697265625, output=0.408216114687
			11'd407: out = 32'b00000000000000000011010001100011; // input=0.39794921875, output=0.409280349921
			11'd408: out = 32'b00000000000000000011010010000110; // input=0.39892578125, output=0.410345076676
			11'd409: out = 32'b00000000000000000011010010101001; // input=0.39990234375, output=0.41141029684
			11'd410: out = 32'b00000000000000000011010011001100; // input=0.40087890625, output=0.412476012313
			11'd411: out = 32'b00000000000000000011010011101111; // input=0.40185546875, output=0.413542224997
			11'd412: out = 32'b00000000000000000011010100010010; // input=0.40283203125, output=0.414608936802
			11'd413: out = 32'b00000000000000000011010100110101; // input=0.40380859375, output=0.415676149646
			11'd414: out = 32'b00000000000000000011010101011000; // input=0.40478515625, output=0.416743865453
			11'd415: out = 32'b00000000000000000011010101111011; // input=0.40576171875, output=0.417812086153
			11'd416: out = 32'b00000000000000000011010110011110; // input=0.40673828125, output=0.418880813684
			11'd417: out = 32'b00000000000000000011010111000001; // input=0.40771484375, output=0.419950049991
			11'd418: out = 32'b00000000000000000011010111100100; // input=0.40869140625, output=0.421019797024
			11'd419: out = 32'b00000000000000000011011000000111; // input=0.40966796875, output=0.422090056743
			11'd420: out = 32'b00000000000000000011011000101010; // input=0.41064453125, output=0.423160831114
			11'd421: out = 32'b00000000000000000011011001001101; // input=0.41162109375, output=0.424232122107
			11'd422: out = 32'b00000000000000000011011001110000; // input=0.41259765625, output=0.425303931704
			11'd423: out = 32'b00000000000000000011011010010011; // input=0.41357421875, output=0.426376261892
			11'd424: out = 32'b00000000000000000011011010110111; // input=0.41455078125, output=0.427449114664
			11'd425: out = 32'b00000000000000000011011011011010; // input=0.41552734375, output=0.428522492022
			11'd426: out = 32'b00000000000000000011011011111101; // input=0.41650390625, output=0.429596395974
			11'd427: out = 32'b00000000000000000011011100100000; // input=0.41748046875, output=0.430670828538
			11'd428: out = 32'b00000000000000000011011101000011; // input=0.41845703125, output=0.431745791736
			11'd429: out = 32'b00000000000000000011011101100111; // input=0.41943359375, output=0.432821287599
			11'd430: out = 32'b00000000000000000011011110001010; // input=0.42041015625, output=0.433897318166
			11'd431: out = 32'b00000000000000000011011110101101; // input=0.42138671875, output=0.434973885483
			11'd432: out = 32'b00000000000000000011011111010001; // input=0.42236328125, output=0.436050991604
			11'd433: out = 32'b00000000000000000011011111110100; // input=0.42333984375, output=0.437128638589
			11'd434: out = 32'b00000000000000000011100000010111; // input=0.42431640625, output=0.438206828509
			11'd435: out = 32'b00000000000000000011100000111011; // input=0.42529296875, output=0.439285563439
			11'd436: out = 32'b00000000000000000011100001011110; // input=0.42626953125, output=0.440364845464
			11'd437: out = 32'b00000000000000000011100010000001; // input=0.42724609375, output=0.441444676676
			11'd438: out = 32'b00000000000000000011100010100101; // input=0.42822265625, output=0.442525059177
			11'd439: out = 32'b00000000000000000011100011001000; // input=0.42919921875, output=0.443605995073
			11'd440: out = 32'b00000000000000000011100011101100; // input=0.43017578125, output=0.444687486481
			11'd441: out = 32'b00000000000000000011100100001111; // input=0.43115234375, output=0.445769535526
			11'd442: out = 32'b00000000000000000011100100110010; // input=0.43212890625, output=0.446852144339
			11'd443: out = 32'b00000000000000000011100101010110; // input=0.43310546875, output=0.447935315062
			11'd444: out = 32'b00000000000000000011100101111001; // input=0.43408203125, output=0.449019049842
			11'd445: out = 32'b00000000000000000011100110011101; // input=0.43505859375, output=0.450103350837
			11'd446: out = 32'b00000000000000000011100111000001; // input=0.43603515625, output=0.451188220212
			11'd447: out = 32'b00000000000000000011100111100100; // input=0.43701171875, output=0.452273660141
			11'd448: out = 32'b00000000000000000011101000001000; // input=0.43798828125, output=0.453359672806
			11'd449: out = 32'b00000000000000000011101000101011; // input=0.43896484375, output=0.454446260396
			11'd450: out = 32'b00000000000000000011101001001111; // input=0.43994140625, output=0.455533425112
			11'd451: out = 32'b00000000000000000011101001110011; // input=0.44091796875, output=0.456621169161
			11'd452: out = 32'b00000000000000000011101010010110; // input=0.44189453125, output=0.457709494758
			11'd453: out = 32'b00000000000000000011101010111010; // input=0.44287109375, output=0.458798404129
			11'd454: out = 32'b00000000000000000011101011011110; // input=0.44384765625, output=0.459887899507
			11'd455: out = 32'b00000000000000000011101100000001; // input=0.44482421875, output=0.460977983136
			11'd456: out = 32'b00000000000000000011101100100101; // input=0.44580078125, output=0.462068657266
			11'd457: out = 32'b00000000000000000011101101001001; // input=0.44677734375, output=0.463159924156
			11'd458: out = 32'b00000000000000000011101101101101; // input=0.44775390625, output=0.464251786078
			11'd459: out = 32'b00000000000000000011101110010000; // input=0.44873046875, output=0.465344245308
			11'd460: out = 32'b00000000000000000011101110110100; // input=0.44970703125, output=0.466437304135
			11'd461: out = 32'b00000000000000000011101111011000; // input=0.45068359375, output=0.467530964854
			11'd462: out = 32'b00000000000000000011101111111100; // input=0.45166015625, output=0.468625229772
			11'd463: out = 32'b00000000000000000011110000100000; // input=0.45263671875, output=0.469720101202
			11'd464: out = 32'b00000000000000000011110001000100; // input=0.45361328125, output=0.47081558147
			11'd465: out = 32'b00000000000000000011110001101000; // input=0.45458984375, output=0.47191167291
			11'd466: out = 32'b00000000000000000011110010001100; // input=0.45556640625, output=0.473008377863
			11'd467: out = 32'b00000000000000000011110010101111; // input=0.45654296875, output=0.474105698684
			11'd468: out = 32'b00000000000000000011110011010011; // input=0.45751953125, output=0.475203637734
			11'd469: out = 32'b00000000000000000011110011110111; // input=0.45849609375, output=0.476302197385
			11'd470: out = 32'b00000000000000000011110100011011; // input=0.45947265625, output=0.477401380019
			11'd471: out = 32'b00000000000000000011110101000000; // input=0.46044921875, output=0.478501188027
			11'd472: out = 32'b00000000000000000011110101100100; // input=0.46142578125, output=0.47960162381
			11'd473: out = 32'b00000000000000000011110110001000; // input=0.46240234375, output=0.48070268978
			11'd474: out = 32'b00000000000000000011110110101100; // input=0.46337890625, output=0.481804388357
			11'd475: out = 32'b00000000000000000011110111010000; // input=0.46435546875, output=0.482906721972
			11'd476: out = 32'b00000000000000000011110111110100; // input=0.46533203125, output=0.484009693068
			11'd477: out = 32'b00000000000000000011111000011000; // input=0.46630859375, output=0.485113304095
			11'd478: out = 32'b00000000000000000011111000111100; // input=0.46728515625, output=0.486217557514
			11'd479: out = 32'b00000000000000000011111001100001; // input=0.46826171875, output=0.487322455798
			11'd480: out = 32'b00000000000000000011111010000101; // input=0.46923828125, output=0.48842800143
			11'd481: out = 32'b00000000000000000011111010101001; // input=0.47021484375, output=0.489534196901
			11'd482: out = 32'b00000000000000000011111011001101; // input=0.47119140625, output=0.490641044716
			11'd483: out = 32'b00000000000000000011111011110010; // input=0.47216796875, output=0.491748547388
			11'd484: out = 32'b00000000000000000011111100010110; // input=0.47314453125, output=0.492856707441
			11'd485: out = 32'b00000000000000000011111100111010; // input=0.47412109375, output=0.493965527411
			11'd486: out = 32'b00000000000000000011111101011111; // input=0.47509765625, output=0.495075009844
			11'd487: out = 32'b00000000000000000011111110000011; // input=0.47607421875, output=0.496185157297
			11'd488: out = 32'b00000000000000000011111110100111; // input=0.47705078125, output=0.497295972337
			11'd489: out = 32'b00000000000000000011111111001100; // input=0.47802734375, output=0.498407457545
			11'd490: out = 32'b00000000000000000011111111110000; // input=0.47900390625, output=0.499519615509
			11'd491: out = 32'b00000000000000000100000000010101; // input=0.47998046875, output=0.500632448832
			11'd492: out = 32'b00000000000000000100000000111001; // input=0.48095703125, output=0.501745960124
			11'd493: out = 32'b00000000000000000100000001011110; // input=0.48193359375, output=0.502860152012
			11'd494: out = 32'b00000000000000000100000010000010; // input=0.48291015625, output=0.503975027128
			11'd495: out = 32'b00000000000000000100000010100111; // input=0.48388671875, output=0.505090588121
			11'd496: out = 32'b00000000000000000100000011001011; // input=0.48486328125, output=0.506206837649
			11'd497: out = 32'b00000000000000000100000011110000; // input=0.48583984375, output=0.50732377838
			11'd498: out = 32'b00000000000000000100000100010101; // input=0.48681640625, output=0.508441412998
			11'd499: out = 32'b00000000000000000100000100111001; // input=0.48779296875, output=0.509559744196
			11'd500: out = 32'b00000000000000000100000101011110; // input=0.48876953125, output=0.510678774679
			11'd501: out = 32'b00000000000000000100000110000011; // input=0.48974609375, output=0.511798507164
			11'd502: out = 32'b00000000000000000100000110100111; // input=0.49072265625, output=0.51291894438
			11'd503: out = 32'b00000000000000000100000111001100; // input=0.49169921875, output=0.51404008907
			11'd504: out = 32'b00000000000000000100000111110001; // input=0.49267578125, output=0.515161943987
			11'd505: out = 32'b00000000000000000100001000010110; // input=0.49365234375, output=0.516284511897
			11'd506: out = 32'b00000000000000000100001000111010; // input=0.49462890625, output=0.517407795578
			11'd507: out = 32'b00000000000000000100001001011111; // input=0.49560546875, output=0.518531797822
			11'd508: out = 32'b00000000000000000100001010000100; // input=0.49658203125, output=0.519656521432
			11'd509: out = 32'b00000000000000000100001010101001; // input=0.49755859375, output=0.520781969224
			11'd510: out = 32'b00000000000000000100001011001110; // input=0.49853515625, output=0.521908144027
			11'd511: out = 32'b00000000000000000100001011110011; // input=0.49951171875, output=0.523035048684
			11'd512: out = 32'b00000000000000000100001100011000; // input=0.50048828125, output=0.524162686048
			11'd513: out = 32'b00000000000000000100001100111101; // input=0.50146484375, output=0.525291058987
			11'd514: out = 32'b00000000000000000100001101100010; // input=0.50244140625, output=0.526420170383
			11'd515: out = 32'b00000000000000000100001110000111; // input=0.50341796875, output=0.527550023129
			11'd516: out = 32'b00000000000000000100001110101100; // input=0.50439453125, output=0.528680620133
			11'd517: out = 32'b00000000000000000100001111010001; // input=0.50537109375, output=0.529811964315
			11'd518: out = 32'b00000000000000000100001111110110; // input=0.50634765625, output=0.53094405861
			11'd519: out = 32'b00000000000000000100010000011011; // input=0.50732421875, output=0.532076905965
			11'd520: out = 32'b00000000000000000100010001000000; // input=0.50830078125, output=0.533210509343
			11'd521: out = 32'b00000000000000000100010001100101; // input=0.50927734375, output=0.534344871718
			11'd522: out = 32'b00000000000000000100010010001011; // input=0.51025390625, output=0.53547999608
			11'd523: out = 32'b00000000000000000100010010110000; // input=0.51123046875, output=0.536615885432
			11'd524: out = 32'b00000000000000000100010011010101; // input=0.51220703125, output=0.537752542791
			11'd525: out = 32'b00000000000000000100010011111010; // input=0.51318359375, output=0.538889971188
			11'd526: out = 32'b00000000000000000100010100100000; // input=0.51416015625, output=0.54002817367
			11'd527: out = 32'b00000000000000000100010101000101; // input=0.51513671875, output=0.541167153296
			11'd528: out = 32'b00000000000000000100010101101010; // input=0.51611328125, output=0.542306913141
			11'd529: out = 32'b00000000000000000100010110010000; // input=0.51708984375, output=0.543447456295
			11'd530: out = 32'b00000000000000000100010110110101; // input=0.51806640625, output=0.544588785861
			11'd531: out = 32'b00000000000000000100010111011011; // input=0.51904296875, output=0.545730904958
			11'd532: out = 32'b00000000000000000100011000000000; // input=0.52001953125, output=0.54687381672
			11'd533: out = 32'b00000000000000000100011000100101; // input=0.52099609375, output=0.548017524295
			11'd534: out = 32'b00000000000000000100011001001011; // input=0.52197265625, output=0.549162030848
			11'd535: out = 32'b00000000000000000100011001110000; // input=0.52294921875, output=0.550307339557
			11'd536: out = 32'b00000000000000000100011010010110; // input=0.52392578125, output=0.551453453618
			11'd537: out = 32'b00000000000000000100011010111100; // input=0.52490234375, output=0.55260037624
			11'd538: out = 32'b00000000000000000100011011100001; // input=0.52587890625, output=0.553748110648
			11'd539: out = 32'b00000000000000000100011100000111; // input=0.52685546875, output=0.554896660084
			11'd540: out = 32'b00000000000000000100011100101101; // input=0.52783203125, output=0.556046027806
			11'd541: out = 32'b00000000000000000100011101010010; // input=0.52880859375, output=0.557196217085
			11'd542: out = 32'b00000000000000000100011101111000; // input=0.52978515625, output=0.558347231212
			11'd543: out = 32'b00000000000000000100011110011110; // input=0.53076171875, output=0.559499073492
			11'd544: out = 32'b00000000000000000100011111000011; // input=0.53173828125, output=0.560651747246
			11'd545: out = 32'b00000000000000000100011111101001; // input=0.53271484375, output=0.561805255813
			11'd546: out = 32'b00000000000000000100100000001111; // input=0.53369140625, output=0.562959602546
			11'd547: out = 32'b00000000000000000100100000110101; // input=0.53466796875, output=0.564114790818
			11'd548: out = 32'b00000000000000000100100001011011; // input=0.53564453125, output=0.565270824016
			11'd549: out = 32'b00000000000000000100100010000001; // input=0.53662109375, output=0.566427705546
			11'd550: out = 32'b00000000000000000100100010100111; // input=0.53759765625, output=0.567585438829
			11'd551: out = 32'b00000000000000000100100011001101; // input=0.53857421875, output=0.568744027306
			11'd552: out = 32'b00000000000000000100100011110011; // input=0.53955078125, output=0.569903474432
			11'd553: out = 32'b00000000000000000100100100011001; // input=0.54052734375, output=0.571063783681
			11'd554: out = 32'b00000000000000000100100100111111; // input=0.54150390625, output=0.572224958546
			11'd555: out = 32'b00000000000000000100100101100101; // input=0.54248046875, output=0.573387002535
			11'd556: out = 32'b00000000000000000100100110001011; // input=0.54345703125, output=0.574549919176
			11'd557: out = 32'b00000000000000000100100110110001; // input=0.54443359375, output=0.575713712013
			11'd558: out = 32'b00000000000000000100100111010111; // input=0.54541015625, output=0.576878384612
			11'd559: out = 32'b00000000000000000100100111111101; // input=0.54638671875, output=0.578043940552
			11'd560: out = 32'b00000000000000000100101000100100; // input=0.54736328125, output=0.579210383434
			11'd561: out = 32'b00000000000000000100101001001010; // input=0.54833984375, output=0.580377716876
			11'd562: out = 32'b00000000000000000100101001110000; // input=0.54931640625, output=0.581545944516
			11'd563: out = 32'b00000000000000000100101010010110; // input=0.55029296875, output=0.58271507001
			11'd564: out = 32'b00000000000000000100101010111101; // input=0.55126953125, output=0.583885097033
			11'd565: out = 32'b00000000000000000100101011100011; // input=0.55224609375, output=0.585056029278
			11'd566: out = 32'b00000000000000000100101100001010; // input=0.55322265625, output=0.586227870461
			11'd567: out = 32'b00000000000000000100101100110000; // input=0.55419921875, output=0.587400624313
			11'd568: out = 32'b00000000000000000100101101010110; // input=0.55517578125, output=0.588574294586
			11'd569: out = 32'b00000000000000000100101101111101; // input=0.55615234375, output=0.589748885055
			11'd570: out = 32'b00000000000000000100101110100011; // input=0.55712890625, output=0.590924399509
			11'd571: out = 32'b00000000000000000100101111001010; // input=0.55810546875, output=0.592100841762
			11'd572: out = 32'b00000000000000000100101111110001; // input=0.55908203125, output=0.593278215646
			11'd573: out = 32'b00000000000000000100110000010111; // input=0.56005859375, output=0.594456525014
			11'd574: out = 32'b00000000000000000100110000111110; // input=0.56103515625, output=0.595635773739
			11'd575: out = 32'b00000000000000000100110001100100; // input=0.56201171875, output=0.596815965716
			11'd576: out = 32'b00000000000000000100110010001011; // input=0.56298828125, output=0.597997104858
			11'd577: out = 32'b00000000000000000100110010110010; // input=0.56396484375, output=0.599179195102
			11'd578: out = 32'b00000000000000000100110011011001; // input=0.56494140625, output=0.600362240405
			11'd579: out = 32'b00000000000000000100110011111111; // input=0.56591796875, output=0.601546244745
			11'd580: out = 32'b00000000000000000100110100100110; // input=0.56689453125, output=0.602731212123
			11'd581: out = 32'b00000000000000000100110101001101; // input=0.56787109375, output=0.60391714656
			11'd582: out = 32'b00000000000000000100110101110100; // input=0.56884765625, output=0.6051040521
			11'd583: out = 32'b00000000000000000100110110011011; // input=0.56982421875, output=0.606291932808
			11'd584: out = 32'b00000000000000000100110111000010; // input=0.57080078125, output=0.607480792772
			11'd585: out = 32'b00000000000000000100110111101001; // input=0.57177734375, output=0.608670636103
			11'd586: out = 32'b00000000000000000100111000010000; // input=0.57275390625, output=0.609861466933
			11'd587: out = 32'b00000000000000000100111000110111; // input=0.57373046875, output=0.611053289418
			11'd588: out = 32'b00000000000000000100111001011110; // input=0.57470703125, output=0.612246107738
			11'd589: out = 32'b00000000000000000100111010000101; // input=0.57568359375, output=0.613439926093
			11'd590: out = 32'b00000000000000000100111010101100; // input=0.57666015625, output=0.614634748708
			11'd591: out = 32'b00000000000000000100111011010100; // input=0.57763671875, output=0.615830579834
			11'd592: out = 32'b00000000000000000100111011111011; // input=0.57861328125, output=0.617027423741
			11'd593: out = 32'b00000000000000000100111100100010; // input=0.57958984375, output=0.618225284727
			11'd594: out = 32'b00000000000000000100111101001001; // input=0.58056640625, output=0.619424167112
			11'd595: out = 32'b00000000000000000100111101110001; // input=0.58154296875, output=0.62062407524
			11'd596: out = 32'b00000000000000000100111110011000; // input=0.58251953125, output=0.621825013482
			11'd597: out = 32'b00000000000000000100111110111111; // input=0.58349609375, output=0.623026986232
			11'd598: out = 32'b00000000000000000100111111100111; // input=0.58447265625, output=0.624229997907
			11'd599: out = 32'b00000000000000000101000000001110; // input=0.58544921875, output=0.625434052954
			11'd600: out = 32'b00000000000000000101000000110110; // input=0.58642578125, output=0.62663915584
			11'd601: out = 32'b00000000000000000101000001011101; // input=0.58740234375, output=0.627845311062
			11'd602: out = 32'b00000000000000000101000010000101; // input=0.58837890625, output=0.629052523141
			11'd603: out = 32'b00000000000000000101000010101100; // input=0.58935546875, output=0.630260796623
			11'd604: out = 32'b00000000000000000101000011010100; // input=0.59033203125, output=0.631470136082
			11'd605: out = 32'b00000000000000000101000011111100; // input=0.59130859375, output=0.632680546116
			11'd606: out = 32'b00000000000000000101000100100011; // input=0.59228515625, output=0.633892031354
			11'd607: out = 32'b00000000000000000101000101001011; // input=0.59326171875, output=0.635104596447
			11'd608: out = 32'b00000000000000000101000101110011; // input=0.59423828125, output=0.636318246077
			11'd609: out = 32'b00000000000000000101000110011011; // input=0.59521484375, output=0.63753298495
			11'd610: out = 32'b00000000000000000101000111000011; // input=0.59619140625, output=0.638748817803
			11'd611: out = 32'b00000000000000000101000111101010; // input=0.59716796875, output=0.639965749399
			11'd612: out = 32'b00000000000000000101001000010010; // input=0.59814453125, output=0.641183784528
			11'd613: out = 32'b00000000000000000101001000111010; // input=0.59912109375, output=0.64240292801
			11'd614: out = 32'b00000000000000000101001001100010; // input=0.60009765625, output=0.643623184695
			11'd615: out = 32'b00000000000000000101001010001010; // input=0.60107421875, output=0.644844559457
			11'd616: out = 32'b00000000000000000101001010110010; // input=0.60205078125, output=0.646067057204
			11'd617: out = 32'b00000000000000000101001011011010; // input=0.60302734375, output=0.647290682871
			11'd618: out = 32'b00000000000000000101001100000011; // input=0.60400390625, output=0.648515441423
			11'd619: out = 32'b00000000000000000101001100101011; // input=0.60498046875, output=0.649741337855
			11'd620: out = 32'b00000000000000000101001101010011; // input=0.60595703125, output=0.650968377191
			11'd621: out = 32'b00000000000000000101001101111011; // input=0.60693359375, output=0.652196564486
			11'd622: out = 32'b00000000000000000101001110100011; // input=0.60791015625, output=0.653425904828
			11'd623: out = 32'b00000000000000000101001111001100; // input=0.60888671875, output=0.654656403331
			11'd624: out = 32'b00000000000000000101001111110100; // input=0.60986328125, output=0.655888065144
			11'd625: out = 32'b00000000000000000101010000011101; // input=0.61083984375, output=0.657120895447
			11'd626: out = 32'b00000000000000000101010001000101; // input=0.61181640625, output=0.658354899451
			11'd627: out = 32'b00000000000000000101010001101101; // input=0.61279296875, output=0.659590082398
			11'd628: out = 32'b00000000000000000101010010010110; // input=0.61376953125, output=0.660826449565
			11'd629: out = 32'b00000000000000000101010010111111; // input=0.61474609375, output=0.662064006259
			11'd630: out = 32'b00000000000000000101010011100111; // input=0.61572265625, output=0.66330275782
			11'd631: out = 32'b00000000000000000101010100010000; // input=0.61669921875, output=0.664542709624
			11'd632: out = 32'b00000000000000000101010100111000; // input=0.61767578125, output=0.665783867077
			11'd633: out = 32'b00000000000000000101010101100001; // input=0.61865234375, output=0.667026235621
			11'd634: out = 32'b00000000000000000101010110001010; // input=0.61962890625, output=0.668269820732
			11'd635: out = 32'b00000000000000000101010110110011; // input=0.62060546875, output=0.669514627918
			11'd636: out = 32'b00000000000000000101010111011011; // input=0.62158203125, output=0.670760662725
			11'd637: out = 32'b00000000000000000101011000000100; // input=0.62255859375, output=0.672007930733
			11'd638: out = 32'b00000000000000000101011000101101; // input=0.62353515625, output=0.673256437555
			11'd639: out = 32'b00000000000000000101011001010110; // input=0.62451171875, output=0.674506188843
			11'd640: out = 32'b00000000000000000101011001111111; // input=0.62548828125, output=0.675757190283
			11'd641: out = 32'b00000000000000000101011010101000; // input=0.62646484375, output=0.677009447598
			11'd642: out = 32'b00000000000000000101011011010001; // input=0.62744140625, output=0.678262966548
			11'd643: out = 32'b00000000000000000101011011111010; // input=0.62841796875, output=0.679517752929
			11'd644: out = 32'b00000000000000000101011100100100; // input=0.62939453125, output=0.680773812575
			11'd645: out = 32'b00000000000000000101011101001101; // input=0.63037109375, output=0.682031151358
			11'd646: out = 32'b00000000000000000101011101110110; // input=0.63134765625, output=0.683289775188
			11'd647: out = 32'b00000000000000000101011110011111; // input=0.63232421875, output=0.684549690012
			11'd648: out = 32'b00000000000000000101011111001001; // input=0.63330078125, output=0.685810901818
			11'd649: out = 32'b00000000000000000101011111110010; // input=0.63427734375, output=0.687073416632
			11'd650: out = 32'b00000000000000000101100000011011; // input=0.63525390625, output=0.688337240519
			11'd651: out = 32'b00000000000000000101100001000101; // input=0.63623046875, output=0.689602379584
			11'd652: out = 32'b00000000000000000101100001101110; // input=0.63720703125, output=0.690868839974
			11'd653: out = 32'b00000000000000000101100010011000; // input=0.63818359375, output=0.692136627875
			11'd654: out = 32'b00000000000000000101100011000010; // input=0.63916015625, output=0.693405749514
			11'd655: out = 32'b00000000000000000101100011101011; // input=0.64013671875, output=0.694676211161
			11'd656: out = 32'b00000000000000000101100100010101; // input=0.64111328125, output=0.695948019125
			11'd657: out = 32'b00000000000000000101100100111111; // input=0.64208984375, output=0.697221179759
			11'd658: out = 32'b00000000000000000101100101101000; // input=0.64306640625, output=0.69849569946
			11'd659: out = 32'b00000000000000000101100110010010; // input=0.64404296875, output=0.699771584666
			11'd660: out = 32'b00000000000000000101100110111100; // input=0.64501953125, output=0.701048841859
			11'd661: out = 32'b00000000000000000101100111100110; // input=0.64599609375, output=0.702327477564
			11'd662: out = 32'b00000000000000000101101000010000; // input=0.64697265625, output=0.703607498353
			11'd663: out = 32'b00000000000000000101101000111010; // input=0.64794921875, output=0.70488891084
			11'd664: out = 32'b00000000000000000101101001100100; // input=0.64892578125, output=0.706171721686
			11'd665: out = 32'b00000000000000000101101010001110; // input=0.64990234375, output=0.707455937596
			11'd666: out = 32'b00000000000000000101101010111000; // input=0.65087890625, output=0.708741565323
			11'd667: out = 32'b00000000000000000101101011100010; // input=0.65185546875, output=0.710028611664
			11'd668: out = 32'b00000000000000000101101100001100; // input=0.65283203125, output=0.711317083466
			11'd669: out = 32'b00000000000000000101101100110111; // input=0.65380859375, output=0.712606987621
			11'd670: out = 32'b00000000000000000101101101100001; // input=0.65478515625, output=0.713898331071
			11'd671: out = 32'b00000000000000000101101110001011; // input=0.65576171875, output=0.715191120804
			11'd672: out = 32'b00000000000000000101101110110110; // input=0.65673828125, output=0.71648536386
			11'd673: out = 32'b00000000000000000101101111100000; // input=0.65771484375, output=0.717781067325
			11'd674: out = 32'b00000000000000000101110000001011; // input=0.65869140625, output=0.719078238338
			11'd675: out = 32'b00000000000000000101110000110101; // input=0.65966796875, output=0.720376884086
			11'd676: out = 32'b00000000000000000101110001100000; // input=0.66064453125, output=0.721677011809
			11'd677: out = 32'b00000000000000000101110010001011; // input=0.66162109375, output=0.722978628796
			11'd678: out = 32'b00000000000000000101110010110101; // input=0.66259765625, output=0.72428174239
			11'd679: out = 32'b00000000000000000101110011100000; // input=0.66357421875, output=0.725586359986
			11'd680: out = 32'b00000000000000000101110100001011; // input=0.66455078125, output=0.726892489032
			11'd681: out = 32'b00000000000000000101110100110110; // input=0.66552734375, output=0.728200137029
			11'd682: out = 32'b00000000000000000101110101100001; // input=0.66650390625, output=0.729509311532
			11'd683: out = 32'b00000000000000000101110110001100; // input=0.66748046875, output=0.730820020153
			11'd684: out = 32'b00000000000000000101110110110111; // input=0.66845703125, output=0.732132270556
			11'd685: out = 32'b00000000000000000101110111100010; // input=0.66943359375, output=0.733446070462
			11'd686: out = 32'b00000000000000000101111000001101; // input=0.67041015625, output=0.734761427651
			11'd687: out = 32'b00000000000000000101111000111000; // input=0.67138671875, output=0.736078349955
			11'd688: out = 32'b00000000000000000101111001100011; // input=0.67236328125, output=0.737396845268
			11'd689: out = 32'b00000000000000000101111010001110; // input=0.67333984375, output=0.73871692154
			11'd690: out = 32'b00000000000000000101111010111010; // input=0.67431640625, output=0.74003858678
			11'd691: out = 32'b00000000000000000101111011100101; // input=0.67529296875, output=0.741361849058
			11'd692: out = 32'b00000000000000000101111100010000; // input=0.67626953125, output=0.742686716502
			11'd693: out = 32'b00000000000000000101111100111100; // input=0.67724609375, output=0.744013197301
			11'd694: out = 32'b00000000000000000101111101100111; // input=0.67822265625, output=0.745341299708
			11'd695: out = 32'b00000000000000000101111110010011; // input=0.67919921875, output=0.746671032034
			11'd696: out = 32'b00000000000000000101111110111111; // input=0.68017578125, output=0.748002402655
			11'd697: out = 32'b00000000000000000101111111101010; // input=0.68115234375, output=0.749335420011
			11'd698: out = 32'b00000000000000000110000000010110; // input=0.68212890625, output=0.750670092604
			11'd699: out = 32'b00000000000000000110000001000010; // input=0.68310546875, output=0.752006429003
			11'd700: out = 32'b00000000000000000110000001101110; // input=0.68408203125, output=0.75334443784
			11'd701: out = 32'b00000000000000000110000010011001; // input=0.68505859375, output=0.754684127815
			11'd702: out = 32'b00000000000000000110000011000101; // input=0.68603515625, output=0.756025507694
			11'd703: out = 32'b00000000000000000110000011110001; // input=0.68701171875, output=0.757368586311
			11'd704: out = 32'b00000000000000000110000100011110; // input=0.68798828125, output=0.758713372569
			11'd705: out = 32'b00000000000000000110000101001010; // input=0.68896484375, output=0.760059875439
			11'd706: out = 32'b00000000000000000110000101110110; // input=0.68994140625, output=0.761408103962
			11'd707: out = 32'b00000000000000000110000110100010; // input=0.69091796875, output=0.76275806725
			11'd708: out = 32'b00000000000000000110000111001110; // input=0.69189453125, output=0.764109774486
			11'd709: out = 32'b00000000000000000110000111111011; // input=0.69287109375, output=0.765463234926
			11'd710: out = 32'b00000000000000000110001000100111; // input=0.69384765625, output=0.766818457899
			11'd711: out = 32'b00000000000000000110001001010100; // input=0.69482421875, output=0.768175452807
			11'd712: out = 32'b00000000000000000110001010000000; // input=0.69580078125, output=0.769534229128
			11'd713: out = 32'b00000000000000000110001010101101; // input=0.69677734375, output=0.770894796414
			11'd714: out = 32'b00000000000000000110001011011001; // input=0.69775390625, output=0.772257164294
			11'd715: out = 32'b00000000000000000110001100000110; // input=0.69873046875, output=0.773621342475
			11'd716: out = 32'b00000000000000000110001100110011; // input=0.69970703125, output=0.774987340742
			11'd717: out = 32'b00000000000000000110001101100000; // input=0.70068359375, output=0.776355168958
			11'd718: out = 32'b00000000000000000110001110001100; // input=0.70166015625, output=0.777724837066
			11'd719: out = 32'b00000000000000000110001110111001; // input=0.70263671875, output=0.779096355093
			11'd720: out = 32'b00000000000000000110001111100110; // input=0.70361328125, output=0.780469733143
			11'd721: out = 32'b00000000000000000110010000010011; // input=0.70458984375, output=0.781844981407
			11'd722: out = 32'b00000000000000000110010001000001; // input=0.70556640625, output=0.783222110157
			11'd723: out = 32'b00000000000000000110010001101110; // input=0.70654296875, output=0.78460112975
			11'd724: out = 32'b00000000000000000110010010011011; // input=0.70751953125, output=0.78598205063
			11'd725: out = 32'b00000000000000000110010011001000; // input=0.70849609375, output=0.787364883328
			11'd726: out = 32'b00000000000000000110010011110110; // input=0.70947265625, output=0.788749638461
			11'd727: out = 32'b00000000000000000110010100100011; // input=0.71044921875, output=0.790136326735
			11'd728: out = 32'b00000000000000000110010101010001; // input=0.71142578125, output=0.791524958947
			11'd729: out = 32'b00000000000000000110010101111110; // input=0.71240234375, output=0.792915545985
			11'd730: out = 32'b00000000000000000110010110101100; // input=0.71337890625, output=0.794308098827
			11'd731: out = 32'b00000000000000000110010111011010; // input=0.71435546875, output=0.795702628547
			11'd732: out = 32'b00000000000000000110011000000111; // input=0.71533203125, output=0.797099146312
			11'd733: out = 32'b00000000000000000110011000110101; // input=0.71630859375, output=0.798497663382
			11'd734: out = 32'b00000000000000000110011001100011; // input=0.71728515625, output=0.799898191117
			11'd735: out = 32'b00000000000000000110011010010001; // input=0.71826171875, output=0.801300740973
			11'd736: out = 32'b00000000000000000110011010111111; // input=0.71923828125, output=0.802705324505
			11'd737: out = 32'b00000000000000000110011011101101; // input=0.72021484375, output=0.804111953369
			11'd738: out = 32'b00000000000000000110011100011011; // input=0.72119140625, output=0.805520639322
			11'd739: out = 32'b00000000000000000110011101001010; // input=0.72216796875, output=0.806931394221
			11'd740: out = 32'b00000000000000000110011101111000; // input=0.72314453125, output=0.808344230032
			11'd741: out = 32'b00000000000000000110011110100110; // input=0.72412109375, output=0.809759158821
			11'd742: out = 32'b00000000000000000110011111010101; // input=0.72509765625, output=0.811176192763
			11'd743: out = 32'b00000000000000000110100000000011; // input=0.72607421875, output=0.812595344141
			11'd744: out = 32'b00000000000000000110100000110010; // input=0.72705078125, output=0.814016625347
			11'd745: out = 32'b00000000000000000110100001100000; // input=0.72802734375, output=0.815440048882
			11'd746: out = 32'b00000000000000000110100010001111; // input=0.72900390625, output=0.816865627361
			11'd747: out = 32'b00000000000000000110100010111110; // input=0.72998046875, output=0.81829337351
			11'd748: out = 32'b00000000000000000110100011101101; // input=0.73095703125, output=0.819723300173
			11'd749: out = 32'b00000000000000000110100100011100; // input=0.73193359375, output=0.821155420307
			11'd750: out = 32'b00000000000000000110100101001011; // input=0.73291015625, output=0.822589746989
			11'd751: out = 32'b00000000000000000110100101111010; // input=0.73388671875, output=0.824026293413
			11'd752: out = 32'b00000000000000000110100110101001; // input=0.73486328125, output=0.825465072897
			11'd753: out = 32'b00000000000000000110100111011000; // input=0.73583984375, output=0.826906098877
			11'd754: out = 32'b00000000000000000110101000000111; // input=0.73681640625, output=0.828349384918
			11'd755: out = 32'b00000000000000000110101000110111; // input=0.73779296875, output=0.829794944707
			11'd756: out = 32'b00000000000000000110101001100110; // input=0.73876953125, output=0.831242792059
			11'd757: out = 32'b00000000000000000110101010010110; // input=0.73974609375, output=0.832692940918
			11'd758: out = 32'b00000000000000000110101011000101; // input=0.74072265625, output=0.834145405359
			11'd759: out = 32'b00000000000000000110101011110101; // input=0.74169921875, output=0.835600199588
			11'd760: out = 32'b00000000000000000110101100100101; // input=0.74267578125, output=0.837057337948
			11'd761: out = 32'b00000000000000000110101101010101; // input=0.74365234375, output=0.838516834915
			11'd762: out = 32'b00000000000000000110101110000100; // input=0.74462890625, output=0.839978705103
			11'd763: out = 32'b00000000000000000110101110110100; // input=0.74560546875, output=0.841442963267
			11'd764: out = 32'b00000000000000000110101111100100; // input=0.74658203125, output=0.842909624303
			11'd765: out = 32'b00000000000000000110110000010101; // input=0.74755859375, output=0.844378703249
			11'd766: out = 32'b00000000000000000110110001000101; // input=0.74853515625, output=0.845850215289
			11'd767: out = 32'b00000000000000000110110001110101; // input=0.74951171875, output=0.847324175756
			11'd768: out = 32'b00000000000000000110110010100101; // input=0.75048828125, output=0.84880060013
			11'd769: out = 32'b00000000000000000110110011010110; // input=0.75146484375, output=0.850279504044
			11'd770: out = 32'b00000000000000000110110100000111; // input=0.75244140625, output=0.851760903282
			11'd771: out = 32'b00000000000000000110110100110111; // input=0.75341796875, output=0.853244813787
			11'd772: out = 32'b00000000000000000110110101101000; // input=0.75439453125, output=0.854731251657
			11'd773: out = 32'b00000000000000000110110110011001; // input=0.75537109375, output=0.856220233152
			11'd774: out = 32'b00000000000000000110110111001001; // input=0.75634765625, output=0.857711774692
			11'd775: out = 32'b00000000000000000110110111111010; // input=0.75732421875, output=0.859205892863
			11'd776: out = 32'b00000000000000000110111000101100; // input=0.75830078125, output=0.860702604419
			11'd777: out = 32'b00000000000000000110111001011101; // input=0.75927734375, output=0.86220192628
			11'd778: out = 32'b00000000000000000110111010001110; // input=0.76025390625, output=0.863703875539
			11'd779: out = 32'b00000000000000000110111010111111; // input=0.76123046875, output=0.865208469465
			11'd780: out = 32'b00000000000000000110111011110001; // input=0.76220703125, output=0.866715725501
			11'd781: out = 32'b00000000000000000110111100100010; // input=0.76318359375, output=0.868225661271
			11'd782: out = 32'b00000000000000000110111101010100; // input=0.76416015625, output=0.869738294579
			11'd783: out = 32'b00000000000000000110111110000101; // input=0.76513671875, output=0.871253643414
			11'd784: out = 32'b00000000000000000110111110110111; // input=0.76611328125, output=0.872771725953
			11'd785: out = 32'b00000000000000000110111111101001; // input=0.76708984375, output=0.874292560562
			11'd786: out = 32'b00000000000000000111000000011011; // input=0.76806640625, output=0.875816165799
			11'd787: out = 32'b00000000000000000111000001001101; // input=0.76904296875, output=0.877342560418
			11'd788: out = 32'b00000000000000000111000001111111; // input=0.77001953125, output=0.878871763373
			11'd789: out = 32'b00000000000000000111000010110001; // input=0.77099609375, output=0.880403793817
			11'd790: out = 32'b00000000000000000111000011100011; // input=0.77197265625, output=0.881938671108
			11'd791: out = 32'b00000000000000000111000100010110; // input=0.77294921875, output=0.883476414811
			11'd792: out = 32'b00000000000000000111000101001000; // input=0.77392578125, output=0.885017044704
			11'd793: out = 32'b00000000000000000111000101111011; // input=0.77490234375, output=0.886560580776
			11'd794: out = 32'b00000000000000000111000110101101; // input=0.77587890625, output=0.888107043235
			11'd795: out = 32'b00000000000000000111000111100000; // input=0.77685546875, output=0.889656452506
			11'd796: out = 32'b00000000000000000111001000010011; // input=0.77783203125, output=0.891208829243
			11'd797: out = 32'b00000000000000000111001001000110; // input=0.77880859375, output=0.892764194322
			11'd798: out = 32'b00000000000000000111001001111001; // input=0.77978515625, output=0.894322568854
			11'd799: out = 32'b00000000000000000111001010101100; // input=0.78076171875, output=0.895883974181
			11'd800: out = 32'b00000000000000000111001011100000; // input=0.78173828125, output=0.897448431885
			11'd801: out = 32'b00000000000000000111001100010011; // input=0.78271484375, output=0.899015963789
			11'd802: out = 32'b00000000000000000111001101000110; // input=0.78369140625, output=0.900586591962
			11'd803: out = 32'b00000000000000000111001101111010; // input=0.78466796875, output=0.902160338722
			11'd804: out = 32'b00000000000000000111001110101110; // input=0.78564453125, output=0.903737226641
			11'd805: out = 32'b00000000000000000111001111100001; // input=0.78662109375, output=0.905317278548
			11'd806: out = 32'b00000000000000000111010000010101; // input=0.78759765625, output=0.906900517533
			11'd807: out = 32'b00000000000000000111010001001001; // input=0.78857421875, output=0.908486966953
			11'd808: out = 32'b00000000000000000111010001111101; // input=0.78955078125, output=0.910076650436
			11'd809: out = 32'b00000000000000000111010010110010; // input=0.79052734375, output=0.911669591883
			11'd810: out = 32'b00000000000000000111010011100110; // input=0.79150390625, output=0.913265815473
			11'd811: out = 32'b00000000000000000111010100011010; // input=0.79248046875, output=0.914865345673
			11'd812: out = 32'b00000000000000000111010101001111; // input=0.79345703125, output=0.916468207233
			11'd813: out = 32'b00000000000000000111010110000011; // input=0.79443359375, output=0.918074425201
			11'd814: out = 32'b00000000000000000111010110111000; // input=0.79541015625, output=0.919684024919
			11'd815: out = 32'b00000000000000000111010111101101; // input=0.79638671875, output=0.921297032036
			11'd816: out = 32'b00000000000000000111011000100010; // input=0.79736328125, output=0.922913472506
			11'd817: out = 32'b00000000000000000111011001010111; // input=0.79833984375, output=0.924533372597
			11'd818: out = 32'b00000000000000000111011010001100; // input=0.79931640625, output=0.926156758898
			11'd819: out = 32'b00000000000000000111011011000010; // input=0.80029296875, output=0.92778365832
			11'd820: out = 32'b00000000000000000111011011110111; // input=0.80126953125, output=0.929414098105
			11'd821: out = 32'b00000000000000000111011100101101; // input=0.80224609375, output=0.931048105828
			11'd822: out = 32'b00000000000000000111011101100010; // input=0.80322265625, output=0.932685709409
			11'd823: out = 32'b00000000000000000111011110011000; // input=0.80419921875, output=0.934326937112
			11'd824: out = 32'b00000000000000000111011111001110; // input=0.80517578125, output=0.935971817557
			11'd825: out = 32'b00000000000000000111100000000100; // input=0.80615234375, output=0.937620379721
			11'd826: out = 32'b00000000000000000111100000111010; // input=0.80712890625, output=0.93927265295
			11'd827: out = 32'b00000000000000000111100001110000; // input=0.80810546875, output=0.940928666959
			11'd828: out = 32'b00000000000000000111100010100111; // input=0.80908203125, output=0.942588451845
			11'd829: out = 32'b00000000000000000111100011011101; // input=0.81005859375, output=0.944252038088
			11'd830: out = 32'b00000000000000000111100100010100; // input=0.81103515625, output=0.945919456565
			11'd831: out = 32'b00000000000000000111100101001011; // input=0.81201171875, output=0.947590738548
			11'd832: out = 32'b00000000000000000111100110000010; // input=0.81298828125, output=0.949265915721
			11'd833: out = 32'b00000000000000000111100110111001; // input=0.81396484375, output=0.95094502018
			11'd834: out = 32'b00000000000000000111100111110000; // input=0.81494140625, output=0.952628084445
			11'd835: out = 32'b00000000000000000111101000100111; // input=0.81591796875, output=0.954315141464
			11'd836: out = 32'b00000000000000000111101001011110; // input=0.81689453125, output=0.956006224626
			11'd837: out = 32'b00000000000000000111101010010110; // input=0.81787109375, output=0.957701367765
			11'd838: out = 32'b00000000000000000111101011001110; // input=0.81884765625, output=0.95940060517
			11'd839: out = 32'b00000000000000000111101100000101; // input=0.81982421875, output=0.961103971595
			11'd840: out = 32'b00000000000000000111101100111101; // input=0.82080078125, output=0.962811502264
			11'd841: out = 32'b00000000000000000111101101110101; // input=0.82177734375, output=0.964523232885
			11'd842: out = 32'b00000000000000000111101110101110; // input=0.82275390625, output=0.966239199654
			11'd843: out = 32'b00000000000000000111101111100110; // input=0.82373046875, output=0.967959439271
			11'd844: out = 32'b00000000000000000111110000011111; // input=0.82470703125, output=0.969683988941
			11'd845: out = 32'b00000000000000000111110001010111; // input=0.82568359375, output=0.971412886393
			11'd846: out = 32'b00000000000000000111110010010000; // input=0.82666015625, output=0.973146169884
			11'd847: out = 32'b00000000000000000111110011001001; // input=0.82763671875, output=0.974883878213
			11'd848: out = 32'b00000000000000000111110100000010; // input=0.82861328125, output=0.976626050731
			11'd849: out = 32'b00000000000000000111110100111011; // input=0.82958984375, output=0.978372727348
			11'd850: out = 32'b00000000000000000111110101110101; // input=0.83056640625, output=0.980123948551
			11'd851: out = 32'b00000000000000000111110110101110; // input=0.83154296875, output=0.981879755413
			11'd852: out = 32'b00000000000000000111110111101000; // input=0.83251953125, output=0.983640189601
			11'd853: out = 32'b00000000000000000111111000100010; // input=0.83349609375, output=0.985405293394
			11'd854: out = 32'b00000000000000000111111001011100; // input=0.83447265625, output=0.987175109694
			11'd855: out = 32'b00000000000000000111111010010110; // input=0.83544921875, output=0.988949682035
			11'd856: out = 32'b00000000000000000111111011010000; // input=0.83642578125, output=0.990729054601
			11'd857: out = 32'b00000000000000000111111100001011; // input=0.83740234375, output=0.992513272239
			11'd858: out = 32'b00000000000000000111111101000101; // input=0.83837890625, output=0.99430238047
			11'd859: out = 32'b00000000000000000111111110000000; // input=0.83935546875, output=0.996096425507
			11'd860: out = 32'b00000000000000000111111110111011; // input=0.84033203125, output=0.997895454266
			11'd861: out = 32'b00000000000000000111111111110110; // input=0.84130859375, output=0.999699514384
			11'd862: out = 32'b00000000000000001000000000110001; // input=0.84228515625, output=1.00150865423
			11'd863: out = 32'b00000000000000001000000001101101; // input=0.84326171875, output=1.00332292294
			11'd864: out = 32'b00000000000000001000000010101001; // input=0.84423828125, output=1.00514237039
			11'd865: out = 32'b00000000000000001000000011100100; // input=0.84521484375, output=1.00696704727
			11'd866: out = 32'b00000000000000001000000100100000; // input=0.84619140625, output=1.00879700506
			11'd867: out = 32'b00000000000000001000000101011100; // input=0.84716796875, output=1.01063229605
			11'd868: out = 32'b00000000000000001000000110011001; // input=0.84814453125, output=1.01247297339
			11'd869: out = 32'b00000000000000001000000111010101; // input=0.84912109375, output=1.01431909107
			11'd870: out = 32'b00000000000000001000001000010010; // input=0.85009765625, output=1.01617070397
			11'd871: out = 32'b00000000000000001000001001001111; // input=0.85107421875, output=1.01802786786
			11'd872: out = 32'b00000000000000001000001010001100; // input=0.85205078125, output=1.01989063942
			11'd873: out = 32'b00000000000000001000001011001001; // input=0.85302734375, output=1.02175907629
			11'd874: out = 32'b00000000000000001000001100000110; // input=0.85400390625, output=1.02363323705
			11'd875: out = 32'b00000000000000001000001101000100; // input=0.85498046875, output=1.02551318129
			11'd876: out = 32'b00000000000000001000001110000010; // input=0.85595703125, output=1.02739896957
			11'd877: out = 32'b00000000000000001000001111000000; // input=0.85693359375, output=1.02929066351
			11'd878: out = 32'b00000000000000001000001111111110; // input=0.85791015625, output=1.03118832579
			11'd879: out = 32'b00000000000000001000010000111100; // input=0.85888671875, output=1.03309202014
			11'd880: out = 32'b00000000000000001000010001111011; // input=0.85986328125, output=1.03500181142
			11'd881: out = 32'b00000000000000001000010010111010; // input=0.86083984375, output=1.03691776563
			11'd882: out = 32'b00000000000000001000010011111001; // input=0.86181640625, output=1.03883994992
			11'd883: out = 32'b00000000000000001000010100111000; // input=0.86279296875, output=1.04076843263
			11'd884: out = 32'b00000000000000001000010101110111; // input=0.86376953125, output=1.04270328333
			11'd885: out = 32'b00000000000000001000010110110111; // input=0.86474609375, output=1.04464457284
			11'd886: out = 32'b00000000000000001000010111110111; // input=0.86572265625, output=1.04659237326
			11'd887: out = 32'b00000000000000001000011000110111; // input=0.86669921875, output=1.04854675801
			11'd888: out = 32'b00000000000000001000011001110111; // input=0.86767578125, output=1.05050780186
			11'd889: out = 32'b00000000000000001000011010111000; // input=0.86865234375, output=1.05247558096
			11'd890: out = 32'b00000000000000001000011011111000; // input=0.86962890625, output=1.0544501729
			11'd891: out = 32'b00000000000000001000011100111001; // input=0.87060546875, output=1.0564316567
			11'd892: out = 32'b00000000000000001000011101111010; // input=0.87158203125, output=1.0584201129
			11'd893: out = 32'b00000000000000001000011110111100; // input=0.87255859375, output=1.06041562356
			11'd894: out = 32'b00000000000000001000011111111101; // input=0.87353515625, output=1.06241827236
			11'd895: out = 32'b00000000000000001000100000111111; // input=0.87451171875, output=1.06442814454
			11'd896: out = 32'b00000000000000001000100010000001; // input=0.87548828125, output=1.06644532706
			11'd897: out = 32'b00000000000000001000100011000100; // input=0.87646484375, output=1.06846990857
			11'd898: out = 32'b00000000000000001000100100000110; // input=0.87744140625, output=1.07050197947
			11'd899: out = 32'b00000000000000001000100101001001; // input=0.87841796875, output=1.07254163199
			11'd900: out = 32'b00000000000000001000100110001100; // input=0.87939453125, output=1.0745889602
			11'd901: out = 32'b00000000000000001000100111001111; // input=0.88037109375, output=1.07664406011
			11'd902: out = 32'b00000000000000001000101000010011; // input=0.88134765625, output=1.07870702967
			11'd903: out = 32'b00000000000000001000101001010111; // input=0.88232421875, output=1.08077796888
			11'd904: out = 32'b00000000000000001000101010011011; // input=0.88330078125, output=1.08285697979
			11'd905: out = 32'b00000000000000001000101011011111; // input=0.88427734375, output=1.08494416663
			11'd906: out = 32'b00000000000000001000101100100100; // input=0.88525390625, output=1.08703963583
			11'd907: out = 32'b00000000000000001000101101101001; // input=0.88623046875, output=1.08914349607
			11'd908: out = 32'b00000000000000001000101110101110; // input=0.88720703125, output=1.09125585841
			11'd909: out = 32'b00000000000000001000101111110100; // input=0.88818359375, output=1.09337683631
			11'd910: out = 32'b00000000000000001000110000111010; // input=0.88916015625, output=1.0955065457
			11'd911: out = 32'b00000000000000001000110010000000; // input=0.89013671875, output=1.0976451051
			11'd912: out = 32'b00000000000000001000110011000110; // input=0.89111328125, output=1.09979263568
			11'd913: out = 32'b00000000000000001000110100001101; // input=0.89208984375, output=1.10194926132
			11'd914: out = 32'b00000000000000001000110101010100; // input=0.89306640625, output=1.10411510871
			11'd915: out = 32'b00000000000000001000110110011011; // input=0.89404296875, output=1.10629030749
			11'd916: out = 32'b00000000000000001000110111100011; // input=0.89501953125, output=1.10847499025
			11'd917: out = 32'b00000000000000001000111000101010; // input=0.89599609375, output=1.1106692927
			11'd918: out = 32'b00000000000000001000111001110011; // input=0.89697265625, output=1.11287335376
			11'd919: out = 32'b00000000000000001000111010111011; // input=0.89794921875, output=1.11508731565
			11'd920: out = 32'b00000000000000001000111100000100; // input=0.89892578125, output=1.117311324
			11'd921: out = 32'b00000000000000001000111101001101; // input=0.89990234375, output=1.11954552799
			11'd922: out = 32'b00000000000000001000111110010111; // input=0.90087890625, output=1.12179008044
			11'd923: out = 32'b00000000000000001000111111100001; // input=0.90185546875, output=1.12404513797
			11'd924: out = 32'b00000000000000001001000000101011; // input=0.90283203125, output=1.1263108611
			11'd925: out = 32'b00000000000000001001000001110110; // input=0.90380859375, output=1.12858741441
			11'd926: out = 32'b00000000000000001001000011000001; // input=0.90478515625, output=1.13087496667
			11'd927: out = 32'b00000000000000001001000100001100; // input=0.90576171875, output=1.13317369102
			11'd928: out = 32'b00000000000000001001000101011000; // input=0.90673828125, output=1.13548376509
			11'd929: out = 32'b00000000000000001001000110100100; // input=0.90771484375, output=1.13780537118
			11'd930: out = 32'b00000000000000001001000111110000; // input=0.90869140625, output=1.14013869645
			11'd931: out = 32'b00000000000000001001001000111101; // input=0.90966796875, output=1.14248393307
			11'd932: out = 32'b00000000000000001001001010001010; // input=0.91064453125, output=1.14484127846
			11'd933: out = 32'b00000000000000001001001011011000; // input=0.91162109375, output=1.14721093543
			11'd934: out = 32'b00000000000000001001001100100110; // input=0.91259765625, output=1.14959311244
			11'd935: out = 32'b00000000000000001001001101110100; // input=0.91357421875, output=1.1519880238
			11'd936: out = 32'b00000000000000001001001111000011; // input=0.91455078125, output=1.1543958899
			11'd937: out = 32'b00000000000000001001010000010011; // input=0.91552734375, output=1.15681693745
			11'd938: out = 32'b00000000000000001001010001100010; // input=0.91650390625, output=1.15925139978
			11'd939: out = 32'b00000000000000001001010010110011; // input=0.91748046875, output=1.16169951703
			11'd940: out = 32'b00000000000000001001010100000011; // input=0.91845703125, output=1.16416153653
			11'd941: out = 32'b00000000000000001001010101010100; // input=0.91943359375, output=1.16663771301
			11'd942: out = 32'b00000000000000001001010110100110; // input=0.92041015625, output=1.16912830899
			11'd943: out = 32'b00000000000000001001010111111000; // input=0.92138671875, output=1.17163359507
			11'd944: out = 32'b00000000000000001001011001001011; // input=0.92236328125, output=1.17415385031
			11'd945: out = 32'b00000000000000001001011010011110; // input=0.92333984375, output=1.17668936258
			11'd946: out = 32'b00000000000000001001011011110001; // input=0.92431640625, output=1.17924042897
			11'd947: out = 32'b00000000000000001001011101000101; // input=0.92529296875, output=1.18180735621
			11'd948: out = 32'b00000000000000001001011110011010; // input=0.92626953125, output=1.1843904611
			11'd949: out = 32'b00000000000000001001011111101111; // input=0.92724609375, output=1.18699007099
			11'd950: out = 32'b00000000000000001001100001000101; // input=0.92822265625, output=1.18960652428
			11'd951: out = 32'b00000000000000001001100010011011; // input=0.92919921875, output=1.19224017094
			11'd952: out = 32'b00000000000000001001100011110010; // input=0.93017578125, output=1.19489137306
			11'd953: out = 32'b00000000000000001001100101001010; // input=0.93115234375, output=1.1975605055
			11'd954: out = 32'b00000000000000001001100110100010; // input=0.93212890625, output=1.20024795643
			11'd955: out = 32'b00000000000000001001100111111010; // input=0.93310546875, output=1.20295412811
			11'd956: out = 32'b00000000000000001001101001010100; // input=0.93408203125, output=1.20567943755
			11'd957: out = 32'b00000000000000001001101010101110; // input=0.93505859375, output=1.20842431728
			11'd958: out = 32'b00000000000000001001101100001000; // input=0.93603515625, output=1.21118921619
			11'd959: out = 32'b00000000000000001001101101100100; // input=0.93701171875, output=1.2139746004
			11'd960: out = 32'b00000000000000001001101110111111; // input=0.93798828125, output=1.21678095422
			11'd961: out = 32'b00000000000000001001110000011100; // input=0.93896484375, output=1.21960878111
			11'd962: out = 32'b00000000000000001001110001111010; // input=0.93994140625, output=1.22245860481
			11'd963: out = 32'b00000000000000001001110011011000; // input=0.94091796875, output=1.22533097047
			11'd964: out = 32'b00000000000000001001110100110111; // input=0.94189453125, output=1.22822644589
			11'd965: out = 32'b00000000000000001001110110010110; // input=0.94287109375, output=1.23114562288
			11'd966: out = 32'b00000000000000001001110111110111; // input=0.94384765625, output=1.23408911871
			11'd967: out = 32'b00000000000000001001111001011000; // input=0.94482421875, output=1.23705757763
			11'd968: out = 32'b00000000000000001001111010111010; // input=0.94580078125, output=1.24005167258
			11'd969: out = 32'b00000000000000001001111100011101; // input=0.94677734375, output=1.24307210702
			11'd970: out = 32'b00000000000000001001111110000001; // input=0.94775390625, output=1.24611961686
			11'd971: out = 32'b00000000000000001001111111100110; // input=0.94873046875, output=1.24919497264
			11'd972: out = 32'b00000000000000001010000001001011; // input=0.94970703125, output=1.25229898181
			11'd973: out = 32'b00000000000000001010000010110010; // input=0.95068359375, output=1.25543249128
			11'd974: out = 32'b00000000000000001010000100011010; // input=0.95166015625, output=1.25859639018
			11'd975: out = 32'b00000000000000001010000110000010; // input=0.95263671875, output=1.26179161284
			11'd976: out = 32'b00000000000000001010000111101100; // input=0.95361328125, output=1.26501914206
			11'd977: out = 32'b00000000000000001010001001010111; // input=0.95458984375, output=1.26828001276
			11'd978: out = 32'b00000000000000001010001011000011; // input=0.95556640625, output=1.27157531586
			11'd979: out = 32'b00000000000000001010001100110000; // input=0.95654296875, output=1.27490620266
			11'd980: out = 32'b00000000000000001010001110011110; // input=0.95751953125, output=1.27827388961
			11'd981: out = 32'b00000000000000001010010000001110; // input=0.95849609375, output=1.28167966359
			11'd982: out = 32'b00000000000000001010010001111111; // input=0.95947265625, output=1.28512488772
			11'd983: out = 32'b00000000000000001010010011110001; // input=0.96044921875, output=1.28861100788
			11'd984: out = 32'b00000000000000001010010101100101; // input=0.96142578125, output=1.2921395599
			11'd985: out = 32'b00000000000000001010010111011010; // input=0.96240234375, output=1.29571217755
			11'd986: out = 32'b00000000000000001010011001010000; // input=0.96337890625, output=1.29933060156
			11'd987: out = 32'b00000000000000001010011011001001; // input=0.96435546875, output=1.30299668967
			11'd988: out = 32'b00000000000000001010011101000010; // input=0.96533203125, output=1.30671242792
			11'd989: out = 32'b00000000000000001010011110111110; // input=0.96630859375, output=1.3104799434
			11'd990: out = 32'b00000000000000001010100000111011; // input=0.96728515625, output=1.31430151869
			11'd991: out = 32'b00000000000000001010100010111010; // input=0.96826171875, output=1.31817960826
			11'd992: out = 32'b00000000000000001010100100111011; // input=0.96923828125, output=1.32211685711
			11'd993: out = 32'b00000000000000001010100110111110; // input=0.97021484375, output=1.32611612215
			11'd994: out = 32'b00000000000000001010101001000011; // input=0.97119140625, output=1.33018049673
			11'd995: out = 32'b00000000000000001010101011001011; // input=0.97216796875, output=1.33431333899
			11'd996: out = 32'b00000000000000001010101101010101; // input=0.97314453125, output=1.33851830468
			11'd997: out = 32'b00000000000000001010101111100001; // input=0.97412109375, output=1.34279938541
			11'd998: out = 32'b00000000000000001010110001110000; // input=0.97509765625, output=1.34716095354
			11'd999: out = 32'b00000000000000001010110100000001; // input=0.97607421875, output=1.35160781497
			11'd1000: out = 32'b00000000000000001010110110010110; // input=0.97705078125, output=1.35614527182
			11'd1001: out = 32'b00000000000000001010111000101110; // input=0.97802734375, output=1.36077919721
			11'd1002: out = 32'b00000000000000001010111011001001; // input=0.97900390625, output=1.36551612523
			11'd1003: out = 32'b00000000000000001010111101101000; // input=0.97998046875, output=1.37036335996
			11'd1004: out = 32'b00000000000000001011000000001011; // input=0.98095703125, output=1.37532910873
			11'd1005: out = 32'b00000000000000001011000010110010; // input=0.98193359375, output=1.38042264672
			11'd1006: out = 32'b00000000000000001011000101011101; // input=0.98291015625, output=1.38565452202
			11'd1007: out = 32'b00000000000000001011001000001101; // input=0.98388671875, output=1.39103681451
			11'd1008: out = 32'b00000000000000001011001011000011; // input=0.98486328125, output=1.39658346647
			11'd1009: out = 32'b00000000000000001011001101111111; // input=0.98583984375, output=1.40231071107
			11'd1010: out = 32'b00000000000000001011010001000001; // input=0.98681640625, output=1.40823763659
			11'd1011: out = 32'b00000000000000001011010100001011; // input=0.98779296875, output=1.41438694293
			11'd1012: out = 32'b00000000000000001011010111011100; // input=0.98876953125, output=1.42078597714
			11'd1013: out = 32'b00000000000000001011011010110111; // input=0.98974609375, output=1.42746818517
			11'd1014: out = 32'b00000000000000001011011110011101; // input=0.99072265625, output=1.43447520447
			11'd1015: out = 32'b00000000000000001011100010001111; // input=0.99169921875, output=1.44185998152
			11'd1016: out = 32'b00000000000000001011100110001111; // input=0.99267578125, output=1.44969160393
			11'd1017: out = 32'b00000000000000001011101010100010; // input=0.99365234375, output=1.45806316311
			11'd1018: out = 32'b00000000000000001011101111001010; // input=0.99462890625, output=1.46710535557
			11'd1019: out = 32'b00000000000000001011110100001111; // input=0.99560546875, output=1.47701196053
			11'd1020: out = 32'b00000000000000001011111001111010; // input=0.99658203125, output=1.48809303047
			11'd1021: out = 32'b00000000000000001100000000011110; // input=0.99755859375, output=1.50090497815
			11'd1022: out = 32'b00000000000000001100001000100010; // input=0.99853515625, output=1.51666312963
			11'd1023: out = 32'b00000000000000001100010100010000; // input=0.99951171875, output=1.53954505509
			11'd1024: out = 32'b10000000000000000000000000010000; // input=-0.00048828125, output=-0.000488281269403
			11'd1025: out = 32'b10000000000000000000000000110000; // input=-0.00146484375, output=-0.00146484427387
			11'd1026: out = 32'b10000000000000000000000001010000; // input=-0.00244140625, output=-0.00244140867533
			11'd1027: out = 32'b10000000000000000000000001110000; // input=-0.00341796875, output=-0.00341797540511
			11'd1028: out = 32'b10000000000000000000000010010000; // input=-0.00439453125, output=-0.00439454539458
			11'd1029: out = 32'b10000000000000000000000010110000; // input=-0.00537109375, output=-0.00537111957513
			11'd1030: out = 32'b10000000000000000000000011010000; // input=-0.00634765625, output=-0.00634769887818
			11'd1031: out = 32'b10000000000000000000000011110000; // input=-0.00732421875, output=-0.0073242842352
			11'd1032: out = 32'b10000000000000000000000100010000; // input=-0.00830078125, output=-0.0083008765777
			11'd1033: out = 32'b10000000000000000000000100110000; // input=-0.00927734375, output=-0.00927747683727
			11'd1034: out = 32'b10000000000000000000000101010000; // input=-0.01025390625, output=-0.0102540859456
			11'd1035: out = 32'b10000000000000000000000101110000; // input=-0.01123046875, output=-0.0112307048343
			11'd1036: out = 32'b10000000000000000000000110010000; // input=-0.01220703125, output=-0.0122073344352
			11'd1037: out = 32'b10000000000000000000000110110000; // input=-0.01318359375, output=-0.0131839756803
			11'd1038: out = 32'b10000000000000000000000111010000; // input=-0.01416015625, output=-0.0141606295016
			11'd1039: out = 32'b10000000000000000000000111110000; // input=-0.01513671875, output=-0.0151372968311
			11'd1040: out = 32'b10000000000000000000001000010000; // input=-0.01611328125, output=-0.016113978601
			11'd1041: out = 32'b10000000000000000000001000110000; // input=-0.01708984375, output=-0.0170906757438
			11'd1042: out = 32'b10000000000000000000001001010000; // input=-0.01806640625, output=-0.0180673891919
			11'd1043: out = 32'b10000000000000000000001001110000; // input=-0.01904296875, output=-0.0190441198779
			11'd1044: out = 32'b10000000000000000000001010010000; // input=-0.02001953125, output=-0.0200208687346
			11'd1045: out = 32'b10000000000000000000001010110000; // input=-0.02099609375, output=-0.0209976366949
			11'd1046: out = 32'b10000000000000000000001011010000; // input=-0.02197265625, output=-0.0219744246919
			11'd1047: out = 32'b10000000000000000000001011110000; // input=-0.02294921875, output=-0.0229512336589
			11'd1048: out = 32'b10000000000000000000001100010000; // input=-0.02392578125, output=-0.0239280645293
			11'd1049: out = 32'b10000000000000000000001100110000; // input=-0.02490234375, output=-0.0249049182366
			11'd1050: out = 32'b10000000000000000000001101010000; // input=-0.02587890625, output=-0.0258817957149
			11'd1051: out = 32'b10000000000000000000001101110000; // input=-0.02685546875, output=-0.026858697898
			11'd1052: out = 32'b10000000000000000000001110010000; // input=-0.02783203125, output=-0.0278356257202
			11'd1053: out = 32'b10000000000000000000001110110000; // input=-0.02880859375, output=-0.028812580116
			11'd1054: out = 32'b10000000000000000000001111010000; // input=-0.02978515625, output=-0.0297895620201
			11'd1055: out = 32'b10000000000000000000001111110000; // input=-0.03076171875, output=-0.0307665723674
			11'd1056: out = 32'b10000000000000000000010000010000; // input=-0.03173828125, output=-0.0317436120931
			11'd1057: out = 32'b10000000000000000000010000110000; // input=-0.03271484375, output=-0.0327206821325
			11'd1058: out = 32'b10000000000000000000010001010000; // input=-0.03369140625, output=-0.0336977834215
			11'd1059: out = 32'b10000000000000000000010001110000; // input=-0.03466796875, output=-0.0346749168959
			11'd1060: out = 32'b10000000000000000000010010010000; // input=-0.03564453125, output=-0.0356520834919
			11'd1061: out = 32'b10000000000000000000010010110000; // input=-0.03662109375, output=-0.0366292841462
			11'd1062: out = 32'b10000000000000000000010011010000; // input=-0.03759765625, output=-0.0376065197954
			11'd1063: out = 32'b10000000000000000000010011110000; // input=-0.03857421875, output=-0.0385837913767
			11'd1064: out = 32'b10000000000000000000010100010000; // input=-0.03955078125, output=-0.0395610998276
			11'd1065: out = 32'b10000000000000000000010100110000; // input=-0.04052734375, output=-0.0405384460857
			11'd1066: out = 32'b10000000000000000000010101010000; // input=-0.04150390625, output=-0.0415158310892
			11'd1067: out = 32'b10000000000000000000010101110000; // input=-0.04248046875, output=-0.0424932557764
			11'd1068: out = 32'b10000000000000000000010110010000; // input=-0.04345703125, output=-0.0434707210861
			11'd1069: out = 32'b10000000000000000000010110110000; // input=-0.04443359375, output=-0.0444482279573
			11'd1070: out = 32'b10000000000000000000010111010001; // input=-0.04541015625, output=-0.0454257773296
			11'd1071: out = 32'b10000000000000000000010111110001; // input=-0.04638671875, output=-0.0464033701426
			11'd1072: out = 32'b10000000000000000000011000010001; // input=-0.04736328125, output=-0.0473810073367
			11'd1073: out = 32'b10000000000000000000011000110001; // input=-0.04833984375, output=-0.0483586898524
			11'd1074: out = 32'b10000000000000000000011001010001; // input=-0.04931640625, output=-0.0493364186307
			11'd1075: out = 32'b10000000000000000000011001110001; // input=-0.05029296875, output=-0.0503141946129
			11'd1076: out = 32'b10000000000000000000011010010001; // input=-0.05126953125, output=-0.0512920187407
			11'd1077: out = 32'b10000000000000000000011010110001; // input=-0.05224609375, output=-0.0522698919565
			11'd1078: out = 32'b10000000000000000000011011010001; // input=-0.05322265625, output=-0.0532478152028
			11'd1079: out = 32'b10000000000000000000011011110001; // input=-0.05419921875, output=-0.0542257894226
			11'd1080: out = 32'b10000000000000000000011100010001; // input=-0.05517578125, output=-0.0552038155595
			11'd1081: out = 32'b10000000000000000000011100110001; // input=-0.05615234375, output=-0.0561818945573
			11'd1082: out = 32'b10000000000000000000011101010001; // input=-0.05712890625, output=-0.0571600273605
			11'd1083: out = 32'b10000000000000000000011101110001; // input=-0.05810546875, output=-0.0581382149139
			11'd1084: out = 32'b10000000000000000000011110010001; // input=-0.05908203125, output=-0.0591164581629
			11'd1085: out = 32'b10000000000000000000011110110001; // input=-0.06005859375, output=-0.0600947580532
			11'd1086: out = 32'b10000000000000000000011111010001; // input=-0.06103515625, output=-0.0610731155313
			11'd1087: out = 32'b10000000000000000000011111110001; // input=-0.06201171875, output=-0.0620515315438
			11'd1088: out = 32'b10000000000000000000100000010001; // input=-0.06298828125, output=-0.0630300070381
			11'd1089: out = 32'b10000000000000000000100000110001; // input=-0.06396484375, output=-0.064008542962
			11'd1090: out = 32'b10000000000000000000100001010001; // input=-0.06494140625, output=-0.064987140264
			11'd1091: out = 32'b10000000000000000000100001110010; // input=-0.06591796875, output=-0.0659657998927
			11'd1092: out = 32'b10000000000000000000100010010010; // input=-0.06689453125, output=-0.0669445227978
			11'd1093: out = 32'b10000000000000000000100010110010; // input=-0.06787109375, output=-0.0679233099292
			11'd1094: out = 32'b10000000000000000000100011010010; // input=-0.06884765625, output=-0.0689021622373
			11'd1095: out = 32'b10000000000000000000100011110010; // input=-0.06982421875, output=-0.0698810806733
			11'd1096: out = 32'b10000000000000000000100100010010; // input=-0.07080078125, output=-0.070860066189
			11'd1097: out = 32'b10000000000000000000100100110010; // input=-0.07177734375, output=-0.0718391197364
			11'd1098: out = 32'b10000000000000000000100101010010; // input=-0.07275390625, output=-0.0728182422686
			11'd1099: out = 32'b10000000000000000000100101110010; // input=-0.07373046875, output=-0.0737974347388
			11'd1100: out = 32'b10000000000000000000100110010010; // input=-0.07470703125, output=-0.0747766981013
			11'd1101: out = 32'b10000000000000000000100110110010; // input=-0.07568359375, output=-0.0757560333106
			11'd1102: out = 32'b10000000000000000000100111010010; // input=-0.07666015625, output=-0.0767354413221
			11'd1103: out = 32'b10000000000000000000100111110011; // input=-0.07763671875, output=-0.0777149230917
			11'd1104: out = 32'b10000000000000000000101000010011; // input=-0.07861328125, output=-0.0786944795761
			11'd1105: out = 32'b10000000000000000000101000110011; // input=-0.07958984375, output=-0.0796741117323
			11'd1106: out = 32'b10000000000000000000101001010011; // input=-0.08056640625, output=-0.0806538205183
			11'd1107: out = 32'b10000000000000000000101001110011; // input=-0.08154296875, output=-0.0816336068927
			11'd1108: out = 32'b10000000000000000000101010010011; // input=-0.08251953125, output=-0.0826134718148
			11'd1109: out = 32'b10000000000000000000101010110011; // input=-0.08349609375, output=-0.0835934162443
			11'd1110: out = 32'b10000000000000000000101011010011; // input=-0.08447265625, output=-0.084573441142
			11'd1111: out = 32'b10000000000000000000101011110011; // input=-0.08544921875, output=-0.0855535474692
			11'd1112: out = 32'b10000000000000000000101100010100; // input=-0.08642578125, output=-0.086533736188
			11'd1113: out = 32'b10000000000000000000101100110100; // input=-0.08740234375, output=-0.087514008261
			11'd1114: out = 32'b10000000000000000000101101010100; // input=-0.08837890625, output=-0.0884943646517
			11'd1115: out = 32'b10000000000000000000101101110100; // input=-0.08935546875, output=-0.0894748063244
			11'd1116: out = 32'b10000000000000000000101110010100; // input=-0.09033203125, output=-0.0904553342441
			11'd1117: out = 32'b10000000000000000000101110110100; // input=-0.09130859375, output=-0.0914359493765
			11'd1118: out = 32'b10000000000000000000101111010100; // input=-0.09228515625, output=-0.0924166526881
			11'd1119: out = 32'b10000000000000000000101111110100; // input=-0.09326171875, output=-0.0933974451461
			11'd1120: out = 32'b10000000000000000000110000010101; // input=-0.09423828125, output=-0.0943783277186
			11'd1121: out = 32'b10000000000000000000110000110101; // input=-0.09521484375, output=-0.0953593013745
			11'd1122: out = 32'b10000000000000000000110001010101; // input=-0.09619140625, output=-0.0963403670833
			11'd1123: out = 32'b10000000000000000000110001110101; // input=-0.09716796875, output=-0.0973215258156
			11'd1124: out = 32'b10000000000000000000110010010101; // input=-0.09814453125, output=-0.0983027785426
			11'd1125: out = 32'b10000000000000000000110010110101; // input=-0.09912109375, output=-0.0992841262364
			11'd1126: out = 32'b10000000000000000000110011010110; // input=-0.10009765625, output=-0.10026556987
			11'd1127: out = 32'b10000000000000000000110011110110; // input=-0.10107421875, output=-0.101247110417
			11'd1128: out = 32'b10000000000000000000110100010110; // input=-0.10205078125, output=-0.102228748852
			11'd1129: out = 32'b10000000000000000000110100110110; // input=-0.10302734375, output=-0.103210486151
			11'd1130: out = 32'b10000000000000000000110101010110; // input=-0.10400390625, output=-0.10419232329
			11'd1131: out = 32'b10000000000000000000110101110110; // input=-0.10498046875, output=-0.105174261246
			11'd1132: out = 32'b10000000000000000000110110010111; // input=-0.10595703125, output=-0.106156300998
			11'd1133: out = 32'b10000000000000000000110110110111; // input=-0.10693359375, output=-0.107138443524
			11'd1134: out = 32'b10000000000000000000110111010111; // input=-0.10791015625, output=-0.108120689804
			11'd1135: out = 32'b10000000000000000000110111110111; // input=-0.10888671875, output=-0.10910304082
			11'd1136: out = 32'b10000000000000000000111000010111; // input=-0.10986328125, output=-0.110085497553
			11'd1137: out = 32'b10000000000000000000111000110111; // input=-0.11083984375, output=-0.111068060986
			11'd1138: out = 32'b10000000000000000000111001011000; // input=-0.11181640625, output=-0.112050732102
			11'd1139: out = 32'b10000000000000000000111001111000; // input=-0.11279296875, output=-0.113033511886
			11'd1140: out = 32'b10000000000000000000111010011000; // input=-0.11376953125, output=-0.114016401324
			11'd1141: out = 32'b10000000000000000000111010111000; // input=-0.11474609375, output=-0.114999401402
			11'd1142: out = 32'b10000000000000000000111011011001; // input=-0.11572265625, output=-0.115982513109
			11'd1143: out = 32'b10000000000000000000111011111001; // input=-0.11669921875, output=-0.116965737431
			11'd1144: out = 32'b10000000000000000000111100011001; // input=-0.11767578125, output=-0.11794907536
			11'd1145: out = 32'b10000000000000000000111100111001; // input=-0.11865234375, output=-0.118932527885
			11'd1146: out = 32'b10000000000000000000111101011001; // input=-0.11962890625, output=-0.119916095998
			11'd1147: out = 32'b10000000000000000000111101111010; // input=-0.12060546875, output=-0.120899780692
			11'd1148: out = 32'b10000000000000000000111110011010; // input=-0.12158203125, output=-0.12188358296
			11'd1149: out = 32'b10000000000000000000111110111010; // input=-0.12255859375, output=-0.122867503798
			11'd1150: out = 32'b10000000000000000000111111011010; // input=-0.12353515625, output=-0.1238515442
			11'd1151: out = 32'b10000000000000000000111111111011; // input=-0.12451171875, output=-0.124835705164
			11'd1152: out = 32'b10000000000000000001000000011011; // input=-0.12548828125, output=-0.125819987687
			11'd1153: out = 32'b10000000000000000001000000111011; // input=-0.12646484375, output=-0.126804392769
			11'd1154: out = 32'b10000000000000000001000001011011; // input=-0.12744140625, output=-0.12778892141
			11'd1155: out = 32'b10000000000000000001000001111100; // input=-0.12841796875, output=-0.12877357461
			11'd1156: out = 32'b10000000000000000001000010011100; // input=-0.12939453125, output=-0.129758353373
			11'd1157: out = 32'b10000000000000000001000010111100; // input=-0.13037109375, output=-0.130743258701
			11'd1158: out = 32'b10000000000000000001000011011100; // input=-0.13134765625, output=-0.1317282916
			11'd1159: out = 32'b10000000000000000001000011111101; // input=-0.13232421875, output=-0.132713453074
			11'd1160: out = 32'b10000000000000000001000100011101; // input=-0.13330078125, output=-0.133698744131
			11'd1161: out = 32'b10000000000000000001000100111101; // input=-0.13427734375, output=-0.134684165779
			11'd1162: out = 32'b10000000000000000001000101011110; // input=-0.13525390625, output=-0.135669719027
			11'd1163: out = 32'b10000000000000000001000101111110; // input=-0.13623046875, output=-0.136655404886
			11'd1164: out = 32'b10000000000000000001000110011110; // input=-0.13720703125, output=-0.137641224367
			11'd1165: out = 32'b10000000000000000001000110111111; // input=-0.13818359375, output=-0.138627178482
			11'd1166: out = 32'b10000000000000000001000111011111; // input=-0.13916015625, output=-0.139613268246
			11'd1167: out = 32'b10000000000000000001000111111111; // input=-0.14013671875, output=-0.140599494675
			11'd1168: out = 32'b10000000000000000001001000011111; // input=-0.14111328125, output=-0.141585858784
			11'd1169: out = 32'b10000000000000000001001001000000; // input=-0.14208984375, output=-0.142572361592
			11'd1170: out = 32'b10000000000000000001001001100000; // input=-0.14306640625, output=-0.143559004117
			11'd1171: out = 32'b10000000000000000001001010000000; // input=-0.14404296875, output=-0.144545787379
			11'd1172: out = 32'b10000000000000000001001010100001; // input=-0.14501953125, output=-0.145532712401
			11'd1173: out = 32'b10000000000000000001001011000001; // input=-0.14599609375, output=-0.146519780204
			11'd1174: out = 32'b10000000000000000001001011100010; // input=-0.14697265625, output=-0.147506991814
			11'd1175: out = 32'b10000000000000000001001100000010; // input=-0.14794921875, output=-0.148494348255
			11'd1176: out = 32'b10000000000000000001001100100010; // input=-0.14892578125, output=-0.149481850554
			11'd1177: out = 32'b10000000000000000001001101000011; // input=-0.14990234375, output=-0.15046949974
			11'd1178: out = 32'b10000000000000000001001101100011; // input=-0.15087890625, output=-0.151457296841
			11'd1179: out = 32'b10000000000000000001001110000011; // input=-0.15185546875, output=-0.152445242889
			11'd1180: out = 32'b10000000000000000001001110100100; // input=-0.15283203125, output=-0.153433338915
			11'd1181: out = 32'b10000000000000000001001111000100; // input=-0.15380859375, output=-0.154421585953
			11'd1182: out = 32'b10000000000000000001001111100100; // input=-0.15478515625, output=-0.155409985038
			11'd1183: out = 32'b10000000000000000001010000000101; // input=-0.15576171875, output=-0.156398537206
			11'd1184: out = 32'b10000000000000000001010000100101; // input=-0.15673828125, output=-0.157387243495
			11'd1185: out = 32'b10000000000000000001010001000110; // input=-0.15771484375, output=-0.158376104944
			11'd1186: out = 32'b10000000000000000001010001100110; // input=-0.15869140625, output=-0.159365122593
			11'd1187: out = 32'b10000000000000000001010010000110; // input=-0.15966796875, output=-0.160354297484
			11'd1188: out = 32'b10000000000000000001010010100111; // input=-0.16064453125, output=-0.161343630661
			11'd1189: out = 32'b10000000000000000001010011000111; // input=-0.16162109375, output=-0.162333123168
			11'd1190: out = 32'b10000000000000000001010011101000; // input=-0.16259765625, output=-0.163322776052
			11'd1191: out = 32'b10000000000000000001010100001000; // input=-0.16357421875, output=-0.16431259036
			11'd1192: out = 32'b10000000000000000001010100101001; // input=-0.16455078125, output=-0.165302567142
			11'd1193: out = 32'b10000000000000000001010101001001; // input=-0.16552734375, output=-0.166292707448
			11'd1194: out = 32'b10000000000000000001010101101010; // input=-0.16650390625, output=-0.167283012331
			11'd1195: out = 32'b10000000000000000001010110001010; // input=-0.16748046875, output=-0.168273482845
			11'd1196: out = 32'b10000000000000000001010110101010; // input=-0.16845703125, output=-0.169264120044
			11'd1197: out = 32'b10000000000000000001010111001011; // input=-0.16943359375, output=-0.170254924986
			11'd1198: out = 32'b10000000000000000001010111101011; // input=-0.17041015625, output=-0.171245898729
			11'd1199: out = 32'b10000000000000000001011000001100; // input=-0.17138671875, output=-0.172237042333
			11'd1200: out = 32'b10000000000000000001011000101100; // input=-0.17236328125, output=-0.173228356859
			11'd1201: out = 32'b10000000000000000001011001001101; // input=-0.17333984375, output=-0.174219843372
			11'd1202: out = 32'b10000000000000000001011001101101; // input=-0.17431640625, output=-0.175211502934
			11'd1203: out = 32'b10000000000000000001011010001110; // input=-0.17529296875, output=-0.176203336613
			11'd1204: out = 32'b10000000000000000001011010101110; // input=-0.17626953125, output=-0.177195345477
			11'd1205: out = 32'b10000000000000000001011011001111; // input=-0.17724609375, output=-0.178187530595
			11'd1206: out = 32'b10000000000000000001011011101111; // input=-0.17822265625, output=-0.179179893039
			11'd1207: out = 32'b10000000000000000001011100010000; // input=-0.17919921875, output=-0.180172433881
			11'd1208: out = 32'b10000000000000000001011100110000; // input=-0.18017578125, output=-0.181165154197
			11'd1209: out = 32'b10000000000000000001011101010001; // input=-0.18115234375, output=-0.182158055061
			11'd1210: out = 32'b10000000000000000001011101110001; // input=-0.18212890625, output=-0.183151137553
			11'd1211: out = 32'b10000000000000000001011110010010; // input=-0.18310546875, output=-0.184144402751
			11'd1212: out = 32'b10000000000000000001011110110011; // input=-0.18408203125, output=-0.185137851738
			11'd1213: out = 32'b10000000000000000001011111010011; // input=-0.18505859375, output=-0.186131485596
			11'd1214: out = 32'b10000000000000000001011111110100; // input=-0.18603515625, output=-0.187125305409
			11'd1215: out = 32'b10000000000000000001100000010100; // input=-0.18701171875, output=-0.188119312266
			11'd1216: out = 32'b10000000000000000001100000110101; // input=-0.18798828125, output=-0.189113507254
			11'd1217: out = 32'b10000000000000000001100001010101; // input=-0.18896484375, output=-0.190107891462
			11'd1218: out = 32'b10000000000000000001100001110110; // input=-0.18994140625, output=-0.191102465984
			11'd1219: out = 32'b10000000000000000001100010010111; // input=-0.19091796875, output=-0.192097231912
			11'd1220: out = 32'b10000000000000000001100010110111; // input=-0.19189453125, output=-0.193092190343
			11'd1221: out = 32'b10000000000000000001100011011000; // input=-0.19287109375, output=-0.194087342373
			11'd1222: out = 32'b10000000000000000001100011111000; // input=-0.19384765625, output=-0.195082689101
			11'd1223: out = 32'b10000000000000000001100100011001; // input=-0.19482421875, output=-0.19607823163
			11'd1224: out = 32'b10000000000000000001100100111010; // input=-0.19580078125, output=-0.19707397106
			11'd1225: out = 32'b10000000000000000001100101011010; // input=-0.19677734375, output=-0.198069908498
			11'd1226: out = 32'b10000000000000000001100101111011; // input=-0.19775390625, output=-0.19906604505
			11'd1227: out = 32'b10000000000000000001100110011100; // input=-0.19873046875, output=-0.200062381825
			11'd1228: out = 32'b10000000000000000001100110111100; // input=-0.19970703125, output=-0.201058919932
			11'd1229: out = 32'b10000000000000000001100111011101; // input=-0.20068359375, output=-0.202055660484
			11'd1230: out = 32'b10000000000000000001100111111110; // input=-0.20166015625, output=-0.203052604596
			11'd1231: out = 32'b10000000000000000001101000011110; // input=-0.20263671875, output=-0.204049753384
			11'd1232: out = 32'b10000000000000000001101000111111; // input=-0.20361328125, output=-0.205047107966
			11'd1233: out = 32'b10000000000000000001101001100000; // input=-0.20458984375, output=-0.206044669461
			11'd1234: out = 32'b10000000000000000001101010000000; // input=-0.20556640625, output=-0.207042438993
			11'd1235: out = 32'b10000000000000000001101010100001; // input=-0.20654296875, output=-0.208040417685
			11'd1236: out = 32'b10000000000000000001101011000010; // input=-0.20751953125, output=-0.209038606664
			11'd1237: out = 32'b10000000000000000001101011100010; // input=-0.20849609375, output=-0.210037007058
			11'd1238: out = 32'b10000000000000000001101100000011; // input=-0.20947265625, output=-0.211035619996
			11'd1239: out = 32'b10000000000000000001101100100100; // input=-0.21044921875, output=-0.212034446612
			11'd1240: out = 32'b10000000000000000001101101000101; // input=-0.21142578125, output=-0.21303348804
			11'd1241: out = 32'b10000000000000000001101101100101; // input=-0.21240234375, output=-0.214032745416
			11'd1242: out = 32'b10000000000000000001101110000110; // input=-0.21337890625, output=-0.215032219878
			11'd1243: out = 32'b10000000000000000001101110100111; // input=-0.21435546875, output=-0.216031912567
			11'd1244: out = 32'b10000000000000000001101111001000; // input=-0.21533203125, output=-0.217031824626
			11'd1245: out = 32'b10000000000000000001101111101000; // input=-0.21630859375, output=-0.218031957201
			11'd1246: out = 32'b10000000000000000001110000001001; // input=-0.21728515625, output=-0.219032311437
			11'd1247: out = 32'b10000000000000000001110000101010; // input=-0.21826171875, output=-0.220032888484
			11'd1248: out = 32'b10000000000000000001110001001011; // input=-0.21923828125, output=-0.221033689493
			11'd1249: out = 32'b10000000000000000001110001101100; // input=-0.22021484375, output=-0.222034715618
			11'd1250: out = 32'b10000000000000000001110010001100; // input=-0.22119140625, output=-0.223035968015
			11'd1251: out = 32'b10000000000000000001110010101101; // input=-0.22216796875, output=-0.224037447841
			11'd1252: out = 32'b10000000000000000001110011001110; // input=-0.22314453125, output=-0.225039156258
			11'd1253: out = 32'b10000000000000000001110011101111; // input=-0.22412109375, output=-0.226041094426
			11'd1254: out = 32'b10000000000000000001110100010000; // input=-0.22509765625, output=-0.227043263512
			11'd1255: out = 32'b10000000000000000001110100110001; // input=-0.22607421875, output=-0.228045664681
			11'd1256: out = 32'b10000000000000000001110101010001; // input=-0.22705078125, output=-0.229048299103
			11'd1257: out = 32'b10000000000000000001110101110010; // input=-0.22802734375, output=-0.23005116795
			11'd1258: out = 32'b10000000000000000001110110010011; // input=-0.22900390625, output=-0.231054272395
			11'd1259: out = 32'b10000000000000000001110110110100; // input=-0.22998046875, output=-0.232057613615
			11'd1260: out = 32'b10000000000000000001110111010101; // input=-0.23095703125, output=-0.233061192788
			11'd1261: out = 32'b10000000000000000001110111110110; // input=-0.23193359375, output=-0.234065011095
			11'd1262: out = 32'b10000000000000000001111000010111; // input=-0.23291015625, output=-0.23506906972
			11'd1263: out = 32'b10000000000000000001111000111000; // input=-0.23388671875, output=-0.236073369847
			11'd1264: out = 32'b10000000000000000001111001011001; // input=-0.23486328125, output=-0.237077912665
			11'd1265: out = 32'b10000000000000000001111001111001; // input=-0.23583984375, output=-0.238082699365
			11'd1266: out = 32'b10000000000000000001111010011010; // input=-0.23681640625, output=-0.239087731139
			11'd1267: out = 32'b10000000000000000001111010111011; // input=-0.23779296875, output=-0.240093009183
			11'd1268: out = 32'b10000000000000000001111011011100; // input=-0.23876953125, output=-0.241098534694
			11'd1269: out = 32'b10000000000000000001111011111101; // input=-0.23974609375, output=-0.242104308872
			11'd1270: out = 32'b10000000000000000001111100011110; // input=-0.24072265625, output=-0.243110332922
			11'd1271: out = 32'b10000000000000000001111100111111; // input=-0.24169921875, output=-0.244116608046
			11'd1272: out = 32'b10000000000000000001111101100000; // input=-0.24267578125, output=-0.245123135455
			11'd1273: out = 32'b10000000000000000001111110000001; // input=-0.24365234375, output=-0.246129916357
			11'd1274: out = 32'b10000000000000000001111110100010; // input=-0.24462890625, output=-0.247136951966
			11'd1275: out = 32'b10000000000000000001111111000011; // input=-0.24560546875, output=-0.248144243497
			11'd1276: out = 32'b10000000000000000001111111100100; // input=-0.24658203125, output=-0.249151792168
			11'd1277: out = 32'b10000000000000000010000000000101; // input=-0.24755859375, output=-0.2501595992
			11'd1278: out = 32'b10000000000000000010000000100110; // input=-0.24853515625, output=-0.251167665816
			11'd1279: out = 32'b10000000000000000010000001000111; // input=-0.24951171875, output=-0.252175993242
			11'd1280: out = 32'b10000000000000000010000001101000; // input=-0.25048828125, output=-0.253184582706
			11'd1281: out = 32'b10000000000000000010000010001001; // input=-0.25146484375, output=-0.25419343544
			11'd1282: out = 32'b10000000000000000010000010101010; // input=-0.25244140625, output=-0.255202552678
			11'd1283: out = 32'b10000000000000000010000011001100; // input=-0.25341796875, output=-0.256211935655
			11'd1284: out = 32'b10000000000000000010000011101101; // input=-0.25439453125, output=-0.257221585612
			11'd1285: out = 32'b10000000000000000010000100001110; // input=-0.25537109375, output=-0.25823150379
			11'd1286: out = 32'b10000000000000000010000100101111; // input=-0.25634765625, output=-0.259241691435
			11'd1287: out = 32'b10000000000000000010000101010000; // input=-0.25732421875, output=-0.260252149793
			11'd1288: out = 32'b10000000000000000010000101110001; // input=-0.25830078125, output=-0.261262880115
			11'd1289: out = 32'b10000000000000000010000110010010; // input=-0.25927734375, output=-0.262273883654
			11'd1290: out = 32'b10000000000000000010000110110011; // input=-0.26025390625, output=-0.263285161666
			11'd1291: out = 32'b10000000000000000010000111010100; // input=-0.26123046875, output=-0.26429671541
			11'd1292: out = 32'b10000000000000000010000111110110; // input=-0.26220703125, output=-0.265308546147
			11'd1293: out = 32'b10000000000000000010001000010111; // input=-0.26318359375, output=-0.266320655141
			11'd1294: out = 32'b10000000000000000010001000111000; // input=-0.26416015625, output=-0.267333043661
			11'd1295: out = 32'b10000000000000000010001001011001; // input=-0.26513671875, output=-0.268345712975
			11'd1296: out = 32'b10000000000000000010001001111010; // input=-0.26611328125, output=-0.269358664358
			11'd1297: out = 32'b10000000000000000010001010011100; // input=-0.26708984375, output=-0.270371899086
			11'd1298: out = 32'b10000000000000000010001010111101; // input=-0.26806640625, output=-0.271385418436
			11'd1299: out = 32'b10000000000000000010001011011110; // input=-0.26904296875, output=-0.272399223693
			11'd1300: out = 32'b10000000000000000010001011111111; // input=-0.27001953125, output=-0.273413316139
			11'd1301: out = 32'b10000000000000000010001100100000; // input=-0.27099609375, output=-0.274427697064
			11'd1302: out = 32'b10000000000000000010001101000010; // input=-0.27197265625, output=-0.275442367758
			11'd1303: out = 32'b10000000000000000010001101100011; // input=-0.27294921875, output=-0.276457329516
			11'd1304: out = 32'b10000000000000000010001110000100; // input=-0.27392578125, output=-0.277472583634
			11'd1305: out = 32'b10000000000000000010001110100101; // input=-0.27490234375, output=-0.278488131412
			11'd1306: out = 32'b10000000000000000010001111000111; // input=-0.27587890625, output=-0.279503974155
			11'd1307: out = 32'b10000000000000000010001111101000; // input=-0.27685546875, output=-0.280520113167
			11'd1308: out = 32'b10000000000000000010010000001001; // input=-0.27783203125, output=-0.28153654976
			11'd1309: out = 32'b10000000000000000010010000101011; // input=-0.27880859375, output=-0.282553285244
			11'd1310: out = 32'b10000000000000000010010001001100; // input=-0.27978515625, output=-0.283570320937
			11'd1311: out = 32'b10000000000000000010010001101101; // input=-0.28076171875, output=-0.284587658157
			11'd1312: out = 32'b10000000000000000010010010001111; // input=-0.28173828125, output=-0.285605298226
			11'd1313: out = 32'b10000000000000000010010010110000; // input=-0.28271484375, output=-0.28662324247
			11'd1314: out = 32'b10000000000000000010010011010001; // input=-0.28369140625, output=-0.287641492218
			11'd1315: out = 32'b10000000000000000010010011110011; // input=-0.28466796875, output=-0.288660048801
			11'd1316: out = 32'b10000000000000000010010100010100; // input=-0.28564453125, output=-0.289678913555
			11'd1317: out = 32'b10000000000000000010010100110110; // input=-0.28662109375, output=-0.290698087817
			11'd1318: out = 32'b10000000000000000010010101010111; // input=-0.28759765625, output=-0.291717572931
			11'd1319: out = 32'b10000000000000000010010101111000; // input=-0.28857421875, output=-0.292737370241
			11'd1320: out = 32'b10000000000000000010010110011010; // input=-0.28955078125, output=-0.293757481095
			11'd1321: out = 32'b10000000000000000010010110111011; // input=-0.29052734375, output=-0.294777906847
			11'd1322: out = 32'b10000000000000000010010111011101; // input=-0.29150390625, output=-0.29579864885
			11'd1323: out = 32'b10000000000000000010010111111110; // input=-0.29248046875, output=-0.296819708463
			11'd1324: out = 32'b10000000000000000010011000100000; // input=-0.29345703125, output=-0.29784108705
			11'd1325: out = 32'b10000000000000000010011001000001; // input=-0.29443359375, output=-0.298862785975
			11'd1326: out = 32'b10000000000000000010011001100011; // input=-0.29541015625, output=-0.299884806608
			11'd1327: out = 32'b10000000000000000010011010000100; // input=-0.29638671875, output=-0.300907150321
			11'd1328: out = 32'b10000000000000000010011010100110; // input=-0.29736328125, output=-0.30192981849
			11'd1329: out = 32'b10000000000000000010011011000111; // input=-0.29833984375, output=-0.302952812495
			11'd1330: out = 32'b10000000000000000010011011101001; // input=-0.29931640625, output=-0.30397613372
			11'd1331: out = 32'b10000000000000000010011100001010; // input=-0.30029296875, output=-0.304999783551
			11'd1332: out = 32'b10000000000000000010011100101100; // input=-0.30126953125, output=-0.306023763378
			11'd1333: out = 32'b10000000000000000010011101001101; // input=-0.30224609375, output=-0.307048074597
			11'd1334: out = 32'b10000000000000000010011101101111; // input=-0.30322265625, output=-0.308072718603
			11'd1335: out = 32'b10000000000000000010011110010001; // input=-0.30419921875, output=-0.309097696799
			11'd1336: out = 32'b10000000000000000010011110110010; // input=-0.30517578125, output=-0.310123010591
			11'd1337: out = 32'b10000000000000000010011111010100; // input=-0.30615234375, output=-0.311148661385
			11'd1338: out = 32'b10000000000000000010011111110101; // input=-0.30712890625, output=-0.312174650596
			11'd1339: out = 32'b10000000000000000010100000010111; // input=-0.30810546875, output=-0.31320097964
			11'd1340: out = 32'b10000000000000000010100000111001; // input=-0.30908203125, output=-0.314227649936
			11'd1341: out = 32'b10000000000000000010100001011010; // input=-0.31005859375, output=-0.315254662909
			11'd1342: out = 32'b10000000000000000010100001111100; // input=-0.31103515625, output=-0.316282019985
			11'd1343: out = 32'b10000000000000000010100010011110; // input=-0.31201171875, output=-0.317309722597
			11'd1344: out = 32'b10000000000000000010100010111111; // input=-0.31298828125, output=-0.318337772181
			11'd1345: out = 32'b10000000000000000010100011100001; // input=-0.31396484375, output=-0.319366170175
			11'd1346: out = 32'b10000000000000000010100100000011; // input=-0.31494140625, output=-0.320394918022
			11'd1347: out = 32'b10000000000000000010100100100100; // input=-0.31591796875, output=-0.32142401717
			11'd1348: out = 32'b10000000000000000010100101000110; // input=-0.31689453125, output=-0.32245346907
			11'd1349: out = 32'b10000000000000000010100101101000; // input=-0.31787109375, output=-0.323483275177
			11'd1350: out = 32'b10000000000000000010100110001010; // input=-0.31884765625, output=-0.32451343695
			11'd1351: out = 32'b10000000000000000010100110101011; // input=-0.31982421875, output=-0.325543955852
			11'd1352: out = 32'b10000000000000000010100111001101; // input=-0.32080078125, output=-0.326574833351
			11'd1353: out = 32'b10000000000000000010100111101111; // input=-0.32177734375, output=-0.327606070917
			11'd1354: out = 32'b10000000000000000010101000010001; // input=-0.32275390625, output=-0.328637670026
			11'd1355: out = 32'b10000000000000000010101000110011; // input=-0.32373046875, output=-0.329669632158
			11'd1356: out = 32'b10000000000000000010101001010100; // input=-0.32470703125, output=-0.330701958797
			11'd1357: out = 32'b10000000000000000010101001110110; // input=-0.32568359375, output=-0.331734651429
			11'd1358: out = 32'b10000000000000000010101010011000; // input=-0.32666015625, output=-0.332767711548
			11'd1359: out = 32'b10000000000000000010101010111010; // input=-0.32763671875, output=-0.333801140649
			11'd1360: out = 32'b10000000000000000010101011011100; // input=-0.32861328125, output=-0.334834940233
			11'd1361: out = 32'b10000000000000000010101011111110; // input=-0.32958984375, output=-0.335869111804
			11'd1362: out = 32'b10000000000000000010101100100000; // input=-0.33056640625, output=-0.336903656873
			11'd1363: out = 32'b10000000000000000010101101000010; // input=-0.33154296875, output=-0.337938576951
			11'd1364: out = 32'b10000000000000000010101101100011; // input=-0.33251953125, output=-0.338973873558
			11'd1365: out = 32'b10000000000000000010101110000101; // input=-0.33349609375, output=-0.340009548215
			11'd1366: out = 32'b10000000000000000010101110100111; // input=-0.33447265625, output=-0.341045602449
			11'd1367: out = 32'b10000000000000000010101111001001; // input=-0.33544921875, output=-0.34208203779
			11'd1368: out = 32'b10000000000000000010101111101011; // input=-0.33642578125, output=-0.343118855775
			11'd1369: out = 32'b10000000000000000010110000001101; // input=-0.33740234375, output=-0.344156057942
			11'd1370: out = 32'b10000000000000000010110000101111; // input=-0.33837890625, output=-0.345193645838
			11'd1371: out = 32'b10000000000000000010110001010001; // input=-0.33935546875, output=-0.346231621009
			11'd1372: out = 32'b10000000000000000010110001110011; // input=-0.34033203125, output=-0.347269985011
			11'd1373: out = 32'b10000000000000000010110010010101; // input=-0.34130859375, output=-0.348308739401
			11'd1374: out = 32'b10000000000000000010110010110111; // input=-0.34228515625, output=-0.349347885742
			11'd1375: out = 32'b10000000000000000010110011011001; // input=-0.34326171875, output=-0.350387425601
			11'd1376: out = 32'b10000000000000000010110011111100; // input=-0.34423828125, output=-0.351427360551
			11'd1377: out = 32'b10000000000000000010110100011110; // input=-0.34521484375, output=-0.352467692167
			11'd1378: out = 32'b10000000000000000010110101000000; // input=-0.34619140625, output=-0.353508422032
			11'd1379: out = 32'b10000000000000000010110101100010; // input=-0.34716796875, output=-0.354549551733
			11'd1380: out = 32'b10000000000000000010110110000100; // input=-0.34814453125, output=-0.355591082858
			11'd1381: out = 32'b10000000000000000010110110100110; // input=-0.34912109375, output=-0.356633017006
			11'd1382: out = 32'b10000000000000000010110111001000; // input=-0.35009765625, output=-0.357675355776
			11'd1383: out = 32'b10000000000000000010110111101010; // input=-0.35107421875, output=-0.358718100774
			11'd1384: out = 32'b10000000000000000010111000001101; // input=-0.35205078125, output=-0.359761253611
			11'd1385: out = 32'b10000000000000000010111000101111; // input=-0.35302734375, output=-0.360804815901
			11'd1386: out = 32'b10000000000000000010111001010001; // input=-0.35400390625, output=-0.361848789265
			11'd1387: out = 32'b10000000000000000010111001110011; // input=-0.35498046875, output=-0.362893175329
			11'd1388: out = 32'b10000000000000000010111010010110; // input=-0.35595703125, output=-0.363937975722
			11'd1389: out = 32'b10000000000000000010111010111000; // input=-0.35693359375, output=-0.364983192081
			11'd1390: out = 32'b10000000000000000010111011011010; // input=-0.35791015625, output=-0.366028826045
			11'd1391: out = 32'b10000000000000000010111011111100; // input=-0.35888671875, output=-0.367074879261
			11'd1392: out = 32'b10000000000000000010111100011111; // input=-0.35986328125, output=-0.368121353378
			11'd1393: out = 32'b10000000000000000010111101000001; // input=-0.36083984375, output=-0.369168250053
			11'd1394: out = 32'b10000000000000000010111101100011; // input=-0.36181640625, output=-0.370215570947
			11'd1395: out = 32'b10000000000000000010111110000110; // input=-0.36279296875, output=-0.371263317726
			11'd1396: out = 32'b10000000000000000010111110101000; // input=-0.36376953125, output=-0.372311492062
			11'd1397: out = 32'b10000000000000000010111111001010; // input=-0.36474609375, output=-0.373360095631
			11'd1398: out = 32'b10000000000000000010111111101101; // input=-0.36572265625, output=-0.374409130116
			11'd1399: out = 32'b10000000000000000011000000001111; // input=-0.36669921875, output=-0.375458597205
			11'd1400: out = 32'b10000000000000000011000000110001; // input=-0.36767578125, output=-0.37650849859
			11'd1401: out = 32'b10000000000000000011000001010100; // input=-0.36865234375, output=-0.377558835969
			11'd1402: out = 32'b10000000000000000011000001110110; // input=-0.36962890625, output=-0.378609611047
			11'd1403: out = 32'b10000000000000000011000010011001; // input=-0.37060546875, output=-0.379660825532
			11'd1404: out = 32'b10000000000000000011000010111011; // input=-0.37158203125, output=-0.38071248114
			11'd1405: out = 32'b10000000000000000011000011011110; // input=-0.37255859375, output=-0.381764579591
			11'd1406: out = 32'b10000000000000000011000100000000; // input=-0.37353515625, output=-0.38281712261
			11'd1407: out = 32'b10000000000000000011000100100011; // input=-0.37451171875, output=-0.38387011193
			11'd1408: out = 32'b10000000000000000011000101000101; // input=-0.37548828125, output=-0.384923549288
			11'd1409: out = 32'b10000000000000000011000101101000; // input=-0.37646484375, output=-0.385977436426
			11'd1410: out = 32'b10000000000000000011000110001010; // input=-0.37744140625, output=-0.387031775094
			11'd1411: out = 32'b10000000000000000011000110101101; // input=-0.37841796875, output=-0.388086567045
			11'd1412: out = 32'b10000000000000000011000111001111; // input=-0.37939453125, output=-0.38914181404
			11'd1413: out = 32'b10000000000000000011000111110010; // input=-0.38037109375, output=-0.390197517845
			11'd1414: out = 32'b10000000000000000011001000010101; // input=-0.38134765625, output=-0.391253680232
			11'd1415: out = 32'b10000000000000000011001000110111; // input=-0.38232421875, output=-0.392310302978
			11'd1416: out = 32'b10000000000000000011001001011010; // input=-0.38330078125, output=-0.393367387867
			11'd1417: out = 32'b10000000000000000011001001111101; // input=-0.38427734375, output=-0.394424936689
			11'd1418: out = 32'b10000000000000000011001010011111; // input=-0.38525390625, output=-0.395482951241
			11'd1419: out = 32'b10000000000000000011001011000010; // input=-0.38623046875, output=-0.396541433322
			11'd1420: out = 32'b10000000000000000011001011100101; // input=-0.38720703125, output=-0.397600384742
			11'd1421: out = 32'b10000000000000000011001100000111; // input=-0.38818359375, output=-0.398659807314
			11'd1422: out = 32'b10000000000000000011001100101010; // input=-0.38916015625, output=-0.399719702858
			11'd1423: out = 32'b10000000000000000011001101001101; // input=-0.39013671875, output=-0.400780073201
			11'd1424: out = 32'b10000000000000000011001101110000; // input=-0.39111328125, output=-0.401840920174
			11'd1425: out = 32'b10000000000000000011001110010010; // input=-0.39208984375, output=-0.402902245618
			11'd1426: out = 32'b10000000000000000011001110110101; // input=-0.39306640625, output=-0.403964051377
			11'd1427: out = 32'b10000000000000000011001111011000; // input=-0.39404296875, output=-0.405026339302
			11'd1428: out = 32'b10000000000000000011001111111011; // input=-0.39501953125, output=-0.406089111252
			11'd1429: out = 32'b10000000000000000011010000011110; // input=-0.39599609375, output=-0.40715236909
			11'd1430: out = 32'b10000000000000000011010001000000; // input=-0.39697265625, output=-0.408216114687
			11'd1431: out = 32'b10000000000000000011010001100011; // input=-0.39794921875, output=-0.409280349921
			11'd1432: out = 32'b10000000000000000011010010000110; // input=-0.39892578125, output=-0.410345076676
			11'd1433: out = 32'b10000000000000000011010010101001; // input=-0.39990234375, output=-0.41141029684
			11'd1434: out = 32'b10000000000000000011010011001100; // input=-0.40087890625, output=-0.412476012313
			11'd1435: out = 32'b10000000000000000011010011101111; // input=-0.40185546875, output=-0.413542224997
			11'd1436: out = 32'b10000000000000000011010100010010; // input=-0.40283203125, output=-0.414608936802
			11'd1437: out = 32'b10000000000000000011010100110101; // input=-0.40380859375, output=-0.415676149646
			11'd1438: out = 32'b10000000000000000011010101011000; // input=-0.40478515625, output=-0.416743865453
			11'd1439: out = 32'b10000000000000000011010101111011; // input=-0.40576171875, output=-0.417812086153
			11'd1440: out = 32'b10000000000000000011010110011110; // input=-0.40673828125, output=-0.418880813684
			11'd1441: out = 32'b10000000000000000011010111000001; // input=-0.40771484375, output=-0.419950049991
			11'd1442: out = 32'b10000000000000000011010111100100; // input=-0.40869140625, output=-0.421019797024
			11'd1443: out = 32'b10000000000000000011011000000111; // input=-0.40966796875, output=-0.422090056743
			11'd1444: out = 32'b10000000000000000011011000101010; // input=-0.41064453125, output=-0.423160831114
			11'd1445: out = 32'b10000000000000000011011001001101; // input=-0.41162109375, output=-0.424232122107
			11'd1446: out = 32'b10000000000000000011011001110000; // input=-0.41259765625, output=-0.425303931704
			11'd1447: out = 32'b10000000000000000011011010010011; // input=-0.41357421875, output=-0.426376261892
			11'd1448: out = 32'b10000000000000000011011010110111; // input=-0.41455078125, output=-0.427449114664
			11'd1449: out = 32'b10000000000000000011011011011010; // input=-0.41552734375, output=-0.428522492022
			11'd1450: out = 32'b10000000000000000011011011111101; // input=-0.41650390625, output=-0.429596395974
			11'd1451: out = 32'b10000000000000000011011100100000; // input=-0.41748046875, output=-0.430670828538
			11'd1452: out = 32'b10000000000000000011011101000011; // input=-0.41845703125, output=-0.431745791736
			11'd1453: out = 32'b10000000000000000011011101100111; // input=-0.41943359375, output=-0.432821287599
			11'd1454: out = 32'b10000000000000000011011110001010; // input=-0.42041015625, output=-0.433897318166
			11'd1455: out = 32'b10000000000000000011011110101101; // input=-0.42138671875, output=-0.434973885483
			11'd1456: out = 32'b10000000000000000011011111010001; // input=-0.42236328125, output=-0.436050991604
			11'd1457: out = 32'b10000000000000000011011111110100; // input=-0.42333984375, output=-0.437128638589
			11'd1458: out = 32'b10000000000000000011100000010111; // input=-0.42431640625, output=-0.438206828509
			11'd1459: out = 32'b10000000000000000011100000111011; // input=-0.42529296875, output=-0.439285563439
			11'd1460: out = 32'b10000000000000000011100001011110; // input=-0.42626953125, output=-0.440364845464
			11'd1461: out = 32'b10000000000000000011100010000001; // input=-0.42724609375, output=-0.441444676676
			11'd1462: out = 32'b10000000000000000011100010100101; // input=-0.42822265625, output=-0.442525059177
			11'd1463: out = 32'b10000000000000000011100011001000; // input=-0.42919921875, output=-0.443605995073
			11'd1464: out = 32'b10000000000000000011100011101100; // input=-0.43017578125, output=-0.444687486481
			11'd1465: out = 32'b10000000000000000011100100001111; // input=-0.43115234375, output=-0.445769535526
			11'd1466: out = 32'b10000000000000000011100100110010; // input=-0.43212890625, output=-0.446852144339
			11'd1467: out = 32'b10000000000000000011100101010110; // input=-0.43310546875, output=-0.447935315062
			11'd1468: out = 32'b10000000000000000011100101111001; // input=-0.43408203125, output=-0.449019049842
			11'd1469: out = 32'b10000000000000000011100110011101; // input=-0.43505859375, output=-0.450103350837
			11'd1470: out = 32'b10000000000000000011100111000001; // input=-0.43603515625, output=-0.451188220212
			11'd1471: out = 32'b10000000000000000011100111100100; // input=-0.43701171875, output=-0.452273660141
			11'd1472: out = 32'b10000000000000000011101000001000; // input=-0.43798828125, output=-0.453359672806
			11'd1473: out = 32'b10000000000000000011101000101011; // input=-0.43896484375, output=-0.454446260396
			11'd1474: out = 32'b10000000000000000011101001001111; // input=-0.43994140625, output=-0.455533425112
			11'd1475: out = 32'b10000000000000000011101001110011; // input=-0.44091796875, output=-0.456621169161
			11'd1476: out = 32'b10000000000000000011101010010110; // input=-0.44189453125, output=-0.457709494758
			11'd1477: out = 32'b10000000000000000011101010111010; // input=-0.44287109375, output=-0.458798404129
			11'd1478: out = 32'b10000000000000000011101011011110; // input=-0.44384765625, output=-0.459887899507
			11'd1479: out = 32'b10000000000000000011101100000001; // input=-0.44482421875, output=-0.460977983136
			11'd1480: out = 32'b10000000000000000011101100100101; // input=-0.44580078125, output=-0.462068657266
			11'd1481: out = 32'b10000000000000000011101101001001; // input=-0.44677734375, output=-0.463159924156
			11'd1482: out = 32'b10000000000000000011101101101101; // input=-0.44775390625, output=-0.464251786078
			11'd1483: out = 32'b10000000000000000011101110010000; // input=-0.44873046875, output=-0.465344245308
			11'd1484: out = 32'b10000000000000000011101110110100; // input=-0.44970703125, output=-0.466437304135
			11'd1485: out = 32'b10000000000000000011101111011000; // input=-0.45068359375, output=-0.467530964854
			11'd1486: out = 32'b10000000000000000011101111111100; // input=-0.45166015625, output=-0.468625229772
			11'd1487: out = 32'b10000000000000000011110000100000; // input=-0.45263671875, output=-0.469720101202
			11'd1488: out = 32'b10000000000000000011110001000100; // input=-0.45361328125, output=-0.47081558147
			11'd1489: out = 32'b10000000000000000011110001101000; // input=-0.45458984375, output=-0.47191167291
			11'd1490: out = 32'b10000000000000000011110010001100; // input=-0.45556640625, output=-0.473008377863
			11'd1491: out = 32'b10000000000000000011110010101111; // input=-0.45654296875, output=-0.474105698684
			11'd1492: out = 32'b10000000000000000011110011010011; // input=-0.45751953125, output=-0.475203637734
			11'd1493: out = 32'b10000000000000000011110011110111; // input=-0.45849609375, output=-0.476302197385
			11'd1494: out = 32'b10000000000000000011110100011011; // input=-0.45947265625, output=-0.477401380019
			11'd1495: out = 32'b10000000000000000011110101000000; // input=-0.46044921875, output=-0.478501188027
			11'd1496: out = 32'b10000000000000000011110101100100; // input=-0.46142578125, output=-0.47960162381
			11'd1497: out = 32'b10000000000000000011110110001000; // input=-0.46240234375, output=-0.48070268978
			11'd1498: out = 32'b10000000000000000011110110101100; // input=-0.46337890625, output=-0.481804388357
			11'd1499: out = 32'b10000000000000000011110111010000; // input=-0.46435546875, output=-0.482906721972
			11'd1500: out = 32'b10000000000000000011110111110100; // input=-0.46533203125, output=-0.484009693068
			11'd1501: out = 32'b10000000000000000011111000011000; // input=-0.46630859375, output=-0.485113304095
			11'd1502: out = 32'b10000000000000000011111000111100; // input=-0.46728515625, output=-0.486217557514
			11'd1503: out = 32'b10000000000000000011111001100001; // input=-0.46826171875, output=-0.487322455798
			11'd1504: out = 32'b10000000000000000011111010000101; // input=-0.46923828125, output=-0.48842800143
			11'd1505: out = 32'b10000000000000000011111010101001; // input=-0.47021484375, output=-0.489534196901
			11'd1506: out = 32'b10000000000000000011111011001101; // input=-0.47119140625, output=-0.490641044716
			11'd1507: out = 32'b10000000000000000011111011110010; // input=-0.47216796875, output=-0.491748547388
			11'd1508: out = 32'b10000000000000000011111100010110; // input=-0.47314453125, output=-0.492856707441
			11'd1509: out = 32'b10000000000000000011111100111010; // input=-0.47412109375, output=-0.493965527411
			11'd1510: out = 32'b10000000000000000011111101011111; // input=-0.47509765625, output=-0.495075009844
			11'd1511: out = 32'b10000000000000000011111110000011; // input=-0.47607421875, output=-0.496185157297
			11'd1512: out = 32'b10000000000000000011111110100111; // input=-0.47705078125, output=-0.497295972337
			11'd1513: out = 32'b10000000000000000011111111001100; // input=-0.47802734375, output=-0.498407457545
			11'd1514: out = 32'b10000000000000000011111111110000; // input=-0.47900390625, output=-0.499519615509
			11'd1515: out = 32'b10000000000000000100000000010101; // input=-0.47998046875, output=-0.500632448832
			11'd1516: out = 32'b10000000000000000100000000111001; // input=-0.48095703125, output=-0.501745960124
			11'd1517: out = 32'b10000000000000000100000001011110; // input=-0.48193359375, output=-0.502860152012
			11'd1518: out = 32'b10000000000000000100000010000010; // input=-0.48291015625, output=-0.503975027128
			11'd1519: out = 32'b10000000000000000100000010100111; // input=-0.48388671875, output=-0.505090588121
			11'd1520: out = 32'b10000000000000000100000011001011; // input=-0.48486328125, output=-0.506206837649
			11'd1521: out = 32'b10000000000000000100000011110000; // input=-0.48583984375, output=-0.50732377838
			11'd1522: out = 32'b10000000000000000100000100010101; // input=-0.48681640625, output=-0.508441412998
			11'd1523: out = 32'b10000000000000000100000100111001; // input=-0.48779296875, output=-0.509559744196
			11'd1524: out = 32'b10000000000000000100000101011110; // input=-0.48876953125, output=-0.510678774679
			11'd1525: out = 32'b10000000000000000100000110000011; // input=-0.48974609375, output=-0.511798507164
			11'd1526: out = 32'b10000000000000000100000110100111; // input=-0.49072265625, output=-0.51291894438
			11'd1527: out = 32'b10000000000000000100000111001100; // input=-0.49169921875, output=-0.51404008907
			11'd1528: out = 32'b10000000000000000100000111110001; // input=-0.49267578125, output=-0.515161943987
			11'd1529: out = 32'b10000000000000000100001000010110; // input=-0.49365234375, output=-0.516284511897
			11'd1530: out = 32'b10000000000000000100001000111010; // input=-0.49462890625, output=-0.517407795578
			11'd1531: out = 32'b10000000000000000100001001011111; // input=-0.49560546875, output=-0.518531797822
			11'd1532: out = 32'b10000000000000000100001010000100; // input=-0.49658203125, output=-0.519656521432
			11'd1533: out = 32'b10000000000000000100001010101001; // input=-0.49755859375, output=-0.520781969224
			11'd1534: out = 32'b10000000000000000100001011001110; // input=-0.49853515625, output=-0.521908144027
			11'd1535: out = 32'b10000000000000000100001011110011; // input=-0.49951171875, output=-0.523035048684
			11'd1536: out = 32'b10000000000000000100001100011000; // input=-0.50048828125, output=-0.524162686048
			11'd1537: out = 32'b10000000000000000100001100111101; // input=-0.50146484375, output=-0.525291058987
			11'd1538: out = 32'b10000000000000000100001101100010; // input=-0.50244140625, output=-0.526420170383
			11'd1539: out = 32'b10000000000000000100001110000111; // input=-0.50341796875, output=-0.527550023129
			11'd1540: out = 32'b10000000000000000100001110101100; // input=-0.50439453125, output=-0.528680620133
			11'd1541: out = 32'b10000000000000000100001111010001; // input=-0.50537109375, output=-0.529811964315
			11'd1542: out = 32'b10000000000000000100001111110110; // input=-0.50634765625, output=-0.53094405861
			11'd1543: out = 32'b10000000000000000100010000011011; // input=-0.50732421875, output=-0.532076905965
			11'd1544: out = 32'b10000000000000000100010001000000; // input=-0.50830078125, output=-0.533210509343
			11'd1545: out = 32'b10000000000000000100010001100101; // input=-0.50927734375, output=-0.534344871718
			11'd1546: out = 32'b10000000000000000100010010001011; // input=-0.51025390625, output=-0.53547999608
			11'd1547: out = 32'b10000000000000000100010010110000; // input=-0.51123046875, output=-0.536615885432
			11'd1548: out = 32'b10000000000000000100010011010101; // input=-0.51220703125, output=-0.537752542791
			11'd1549: out = 32'b10000000000000000100010011111010; // input=-0.51318359375, output=-0.538889971188
			11'd1550: out = 32'b10000000000000000100010100100000; // input=-0.51416015625, output=-0.54002817367
			11'd1551: out = 32'b10000000000000000100010101000101; // input=-0.51513671875, output=-0.541167153296
			11'd1552: out = 32'b10000000000000000100010101101010; // input=-0.51611328125, output=-0.542306913141
			11'd1553: out = 32'b10000000000000000100010110010000; // input=-0.51708984375, output=-0.543447456295
			11'd1554: out = 32'b10000000000000000100010110110101; // input=-0.51806640625, output=-0.544588785861
			11'd1555: out = 32'b10000000000000000100010111011011; // input=-0.51904296875, output=-0.545730904958
			11'd1556: out = 32'b10000000000000000100011000000000; // input=-0.52001953125, output=-0.54687381672
			11'd1557: out = 32'b10000000000000000100011000100101; // input=-0.52099609375, output=-0.548017524295
			11'd1558: out = 32'b10000000000000000100011001001011; // input=-0.52197265625, output=-0.549162030848
			11'd1559: out = 32'b10000000000000000100011001110000; // input=-0.52294921875, output=-0.550307339557
			11'd1560: out = 32'b10000000000000000100011010010110; // input=-0.52392578125, output=-0.551453453618
			11'd1561: out = 32'b10000000000000000100011010111100; // input=-0.52490234375, output=-0.55260037624
			11'd1562: out = 32'b10000000000000000100011011100001; // input=-0.52587890625, output=-0.553748110648
			11'd1563: out = 32'b10000000000000000100011100000111; // input=-0.52685546875, output=-0.554896660084
			11'd1564: out = 32'b10000000000000000100011100101101; // input=-0.52783203125, output=-0.556046027806
			11'd1565: out = 32'b10000000000000000100011101010010; // input=-0.52880859375, output=-0.557196217085
			11'd1566: out = 32'b10000000000000000100011101111000; // input=-0.52978515625, output=-0.558347231212
			11'd1567: out = 32'b10000000000000000100011110011110; // input=-0.53076171875, output=-0.559499073492
			11'd1568: out = 32'b10000000000000000100011111000011; // input=-0.53173828125, output=-0.560651747246
			11'd1569: out = 32'b10000000000000000100011111101001; // input=-0.53271484375, output=-0.561805255813
			11'd1570: out = 32'b10000000000000000100100000001111; // input=-0.53369140625, output=-0.562959602546
			11'd1571: out = 32'b10000000000000000100100000110101; // input=-0.53466796875, output=-0.564114790818
			11'd1572: out = 32'b10000000000000000100100001011011; // input=-0.53564453125, output=-0.565270824016
			11'd1573: out = 32'b10000000000000000100100010000001; // input=-0.53662109375, output=-0.566427705546
			11'd1574: out = 32'b10000000000000000100100010100111; // input=-0.53759765625, output=-0.567585438829
			11'd1575: out = 32'b10000000000000000100100011001101; // input=-0.53857421875, output=-0.568744027306
			11'd1576: out = 32'b10000000000000000100100011110011; // input=-0.53955078125, output=-0.569903474432
			11'd1577: out = 32'b10000000000000000100100100011001; // input=-0.54052734375, output=-0.571063783681
			11'd1578: out = 32'b10000000000000000100100100111111; // input=-0.54150390625, output=-0.572224958546
			11'd1579: out = 32'b10000000000000000100100101100101; // input=-0.54248046875, output=-0.573387002535
			11'd1580: out = 32'b10000000000000000100100110001011; // input=-0.54345703125, output=-0.574549919176
			11'd1581: out = 32'b10000000000000000100100110110001; // input=-0.54443359375, output=-0.575713712013
			11'd1582: out = 32'b10000000000000000100100111010111; // input=-0.54541015625, output=-0.576878384612
			11'd1583: out = 32'b10000000000000000100100111111101; // input=-0.54638671875, output=-0.578043940552
			11'd1584: out = 32'b10000000000000000100101000100100; // input=-0.54736328125, output=-0.579210383434
			11'd1585: out = 32'b10000000000000000100101001001010; // input=-0.54833984375, output=-0.580377716876
			11'd1586: out = 32'b10000000000000000100101001110000; // input=-0.54931640625, output=-0.581545944516
			11'd1587: out = 32'b10000000000000000100101010010110; // input=-0.55029296875, output=-0.58271507001
			11'd1588: out = 32'b10000000000000000100101010111101; // input=-0.55126953125, output=-0.583885097033
			11'd1589: out = 32'b10000000000000000100101011100011; // input=-0.55224609375, output=-0.585056029278
			11'd1590: out = 32'b10000000000000000100101100001010; // input=-0.55322265625, output=-0.586227870461
			11'd1591: out = 32'b10000000000000000100101100110000; // input=-0.55419921875, output=-0.587400624313
			11'd1592: out = 32'b10000000000000000100101101010110; // input=-0.55517578125, output=-0.588574294586
			11'd1593: out = 32'b10000000000000000100101101111101; // input=-0.55615234375, output=-0.589748885055
			11'd1594: out = 32'b10000000000000000100101110100011; // input=-0.55712890625, output=-0.590924399509
			11'd1595: out = 32'b10000000000000000100101111001010; // input=-0.55810546875, output=-0.592100841762
			11'd1596: out = 32'b10000000000000000100101111110001; // input=-0.55908203125, output=-0.593278215646
			11'd1597: out = 32'b10000000000000000100110000010111; // input=-0.56005859375, output=-0.594456525014
			11'd1598: out = 32'b10000000000000000100110000111110; // input=-0.56103515625, output=-0.595635773739
			11'd1599: out = 32'b10000000000000000100110001100100; // input=-0.56201171875, output=-0.596815965716
			11'd1600: out = 32'b10000000000000000100110010001011; // input=-0.56298828125, output=-0.597997104858
			11'd1601: out = 32'b10000000000000000100110010110010; // input=-0.56396484375, output=-0.599179195102
			11'd1602: out = 32'b10000000000000000100110011011001; // input=-0.56494140625, output=-0.600362240405
			11'd1603: out = 32'b10000000000000000100110011111111; // input=-0.56591796875, output=-0.601546244745
			11'd1604: out = 32'b10000000000000000100110100100110; // input=-0.56689453125, output=-0.602731212123
			11'd1605: out = 32'b10000000000000000100110101001101; // input=-0.56787109375, output=-0.60391714656
			11'd1606: out = 32'b10000000000000000100110101110100; // input=-0.56884765625, output=-0.6051040521
			11'd1607: out = 32'b10000000000000000100110110011011; // input=-0.56982421875, output=-0.606291932808
			11'd1608: out = 32'b10000000000000000100110111000010; // input=-0.57080078125, output=-0.607480792772
			11'd1609: out = 32'b10000000000000000100110111101001; // input=-0.57177734375, output=-0.608670636103
			11'd1610: out = 32'b10000000000000000100111000010000; // input=-0.57275390625, output=-0.609861466933
			11'd1611: out = 32'b10000000000000000100111000110111; // input=-0.57373046875, output=-0.611053289418
			11'd1612: out = 32'b10000000000000000100111001011110; // input=-0.57470703125, output=-0.612246107738
			11'd1613: out = 32'b10000000000000000100111010000101; // input=-0.57568359375, output=-0.613439926093
			11'd1614: out = 32'b10000000000000000100111010101100; // input=-0.57666015625, output=-0.614634748708
			11'd1615: out = 32'b10000000000000000100111011010100; // input=-0.57763671875, output=-0.615830579834
			11'd1616: out = 32'b10000000000000000100111011111011; // input=-0.57861328125, output=-0.617027423741
			11'd1617: out = 32'b10000000000000000100111100100010; // input=-0.57958984375, output=-0.618225284727
			11'd1618: out = 32'b10000000000000000100111101001001; // input=-0.58056640625, output=-0.619424167112
			11'd1619: out = 32'b10000000000000000100111101110001; // input=-0.58154296875, output=-0.62062407524
			11'd1620: out = 32'b10000000000000000100111110011000; // input=-0.58251953125, output=-0.621825013482
			11'd1621: out = 32'b10000000000000000100111110111111; // input=-0.58349609375, output=-0.623026986232
			11'd1622: out = 32'b10000000000000000100111111100111; // input=-0.58447265625, output=-0.624229997907
			11'd1623: out = 32'b10000000000000000101000000001110; // input=-0.58544921875, output=-0.625434052954
			11'd1624: out = 32'b10000000000000000101000000110110; // input=-0.58642578125, output=-0.62663915584
			11'd1625: out = 32'b10000000000000000101000001011101; // input=-0.58740234375, output=-0.627845311062
			11'd1626: out = 32'b10000000000000000101000010000101; // input=-0.58837890625, output=-0.629052523141
			11'd1627: out = 32'b10000000000000000101000010101100; // input=-0.58935546875, output=-0.630260796623
			11'd1628: out = 32'b10000000000000000101000011010100; // input=-0.59033203125, output=-0.631470136082
			11'd1629: out = 32'b10000000000000000101000011111100; // input=-0.59130859375, output=-0.632680546116
			11'd1630: out = 32'b10000000000000000101000100100011; // input=-0.59228515625, output=-0.633892031354
			11'd1631: out = 32'b10000000000000000101000101001011; // input=-0.59326171875, output=-0.635104596447
			11'd1632: out = 32'b10000000000000000101000101110011; // input=-0.59423828125, output=-0.636318246077
			11'd1633: out = 32'b10000000000000000101000110011011; // input=-0.59521484375, output=-0.63753298495
			11'd1634: out = 32'b10000000000000000101000111000011; // input=-0.59619140625, output=-0.638748817803
			11'd1635: out = 32'b10000000000000000101000111101010; // input=-0.59716796875, output=-0.639965749399
			11'd1636: out = 32'b10000000000000000101001000010010; // input=-0.59814453125, output=-0.641183784528
			11'd1637: out = 32'b10000000000000000101001000111010; // input=-0.59912109375, output=-0.64240292801
			11'd1638: out = 32'b10000000000000000101001001100010; // input=-0.60009765625, output=-0.643623184695
			11'd1639: out = 32'b10000000000000000101001010001010; // input=-0.60107421875, output=-0.644844559457
			11'd1640: out = 32'b10000000000000000101001010110010; // input=-0.60205078125, output=-0.646067057204
			11'd1641: out = 32'b10000000000000000101001011011010; // input=-0.60302734375, output=-0.647290682871
			11'd1642: out = 32'b10000000000000000101001100000011; // input=-0.60400390625, output=-0.648515441423
			11'd1643: out = 32'b10000000000000000101001100101011; // input=-0.60498046875, output=-0.649741337855
			11'd1644: out = 32'b10000000000000000101001101010011; // input=-0.60595703125, output=-0.650968377191
			11'd1645: out = 32'b10000000000000000101001101111011; // input=-0.60693359375, output=-0.652196564486
			11'd1646: out = 32'b10000000000000000101001110100011; // input=-0.60791015625, output=-0.653425904828
			11'd1647: out = 32'b10000000000000000101001111001100; // input=-0.60888671875, output=-0.654656403331
			11'd1648: out = 32'b10000000000000000101001111110100; // input=-0.60986328125, output=-0.655888065144
			11'd1649: out = 32'b10000000000000000101010000011101; // input=-0.61083984375, output=-0.657120895447
			11'd1650: out = 32'b10000000000000000101010001000101; // input=-0.61181640625, output=-0.658354899451
			11'd1651: out = 32'b10000000000000000101010001101101; // input=-0.61279296875, output=-0.659590082398
			11'd1652: out = 32'b10000000000000000101010010010110; // input=-0.61376953125, output=-0.660826449565
			11'd1653: out = 32'b10000000000000000101010010111111; // input=-0.61474609375, output=-0.662064006259
			11'd1654: out = 32'b10000000000000000101010011100111; // input=-0.61572265625, output=-0.66330275782
			11'd1655: out = 32'b10000000000000000101010100010000; // input=-0.61669921875, output=-0.664542709624
			11'd1656: out = 32'b10000000000000000101010100111000; // input=-0.61767578125, output=-0.665783867077
			11'd1657: out = 32'b10000000000000000101010101100001; // input=-0.61865234375, output=-0.667026235621
			11'd1658: out = 32'b10000000000000000101010110001010; // input=-0.61962890625, output=-0.668269820732
			11'd1659: out = 32'b10000000000000000101010110110011; // input=-0.62060546875, output=-0.669514627918
			11'd1660: out = 32'b10000000000000000101010111011011; // input=-0.62158203125, output=-0.670760662725
			11'd1661: out = 32'b10000000000000000101011000000100; // input=-0.62255859375, output=-0.672007930733
			11'd1662: out = 32'b10000000000000000101011000101101; // input=-0.62353515625, output=-0.673256437555
			11'd1663: out = 32'b10000000000000000101011001010110; // input=-0.62451171875, output=-0.674506188843
			11'd1664: out = 32'b10000000000000000101011001111111; // input=-0.62548828125, output=-0.675757190283
			11'd1665: out = 32'b10000000000000000101011010101000; // input=-0.62646484375, output=-0.677009447598
			11'd1666: out = 32'b10000000000000000101011011010001; // input=-0.62744140625, output=-0.678262966548
			11'd1667: out = 32'b10000000000000000101011011111010; // input=-0.62841796875, output=-0.679517752929
			11'd1668: out = 32'b10000000000000000101011100100100; // input=-0.62939453125, output=-0.680773812575
			11'd1669: out = 32'b10000000000000000101011101001101; // input=-0.63037109375, output=-0.682031151358
			11'd1670: out = 32'b10000000000000000101011101110110; // input=-0.63134765625, output=-0.683289775188
			11'd1671: out = 32'b10000000000000000101011110011111; // input=-0.63232421875, output=-0.684549690012
			11'd1672: out = 32'b10000000000000000101011111001001; // input=-0.63330078125, output=-0.685810901818
			11'd1673: out = 32'b10000000000000000101011111110010; // input=-0.63427734375, output=-0.687073416632
			11'd1674: out = 32'b10000000000000000101100000011011; // input=-0.63525390625, output=-0.688337240519
			11'd1675: out = 32'b10000000000000000101100001000101; // input=-0.63623046875, output=-0.689602379584
			11'd1676: out = 32'b10000000000000000101100001101110; // input=-0.63720703125, output=-0.690868839974
			11'd1677: out = 32'b10000000000000000101100010011000; // input=-0.63818359375, output=-0.692136627875
			11'd1678: out = 32'b10000000000000000101100011000010; // input=-0.63916015625, output=-0.693405749514
			11'd1679: out = 32'b10000000000000000101100011101011; // input=-0.64013671875, output=-0.694676211161
			11'd1680: out = 32'b10000000000000000101100100010101; // input=-0.64111328125, output=-0.695948019125
			11'd1681: out = 32'b10000000000000000101100100111111; // input=-0.64208984375, output=-0.697221179759
			11'd1682: out = 32'b10000000000000000101100101101000; // input=-0.64306640625, output=-0.69849569946
			11'd1683: out = 32'b10000000000000000101100110010010; // input=-0.64404296875, output=-0.699771584666
			11'd1684: out = 32'b10000000000000000101100110111100; // input=-0.64501953125, output=-0.701048841859
			11'd1685: out = 32'b10000000000000000101100111100110; // input=-0.64599609375, output=-0.702327477564
			11'd1686: out = 32'b10000000000000000101101000010000; // input=-0.64697265625, output=-0.703607498353
			11'd1687: out = 32'b10000000000000000101101000111010; // input=-0.64794921875, output=-0.70488891084
			11'd1688: out = 32'b10000000000000000101101001100100; // input=-0.64892578125, output=-0.706171721686
			11'd1689: out = 32'b10000000000000000101101010001110; // input=-0.64990234375, output=-0.707455937596
			11'd1690: out = 32'b10000000000000000101101010111000; // input=-0.65087890625, output=-0.708741565323
			11'd1691: out = 32'b10000000000000000101101011100010; // input=-0.65185546875, output=-0.710028611664
			11'd1692: out = 32'b10000000000000000101101100001100; // input=-0.65283203125, output=-0.711317083466
			11'd1693: out = 32'b10000000000000000101101100110111; // input=-0.65380859375, output=-0.712606987621
			11'd1694: out = 32'b10000000000000000101101101100001; // input=-0.65478515625, output=-0.713898331071
			11'd1695: out = 32'b10000000000000000101101110001011; // input=-0.65576171875, output=-0.715191120804
			11'd1696: out = 32'b10000000000000000101101110110110; // input=-0.65673828125, output=-0.71648536386
			11'd1697: out = 32'b10000000000000000101101111100000; // input=-0.65771484375, output=-0.717781067325
			11'd1698: out = 32'b10000000000000000101110000001011; // input=-0.65869140625, output=-0.719078238338
			11'd1699: out = 32'b10000000000000000101110000110101; // input=-0.65966796875, output=-0.720376884086
			11'd1700: out = 32'b10000000000000000101110001100000; // input=-0.66064453125, output=-0.721677011809
			11'd1701: out = 32'b10000000000000000101110010001011; // input=-0.66162109375, output=-0.722978628796
			11'd1702: out = 32'b10000000000000000101110010110101; // input=-0.66259765625, output=-0.72428174239
			11'd1703: out = 32'b10000000000000000101110011100000; // input=-0.66357421875, output=-0.725586359986
			11'd1704: out = 32'b10000000000000000101110100001011; // input=-0.66455078125, output=-0.726892489032
			11'd1705: out = 32'b10000000000000000101110100110110; // input=-0.66552734375, output=-0.728200137029
			11'd1706: out = 32'b10000000000000000101110101100001; // input=-0.66650390625, output=-0.729509311532
			11'd1707: out = 32'b10000000000000000101110110001100; // input=-0.66748046875, output=-0.730820020153
			11'd1708: out = 32'b10000000000000000101110110110111; // input=-0.66845703125, output=-0.732132270556
			11'd1709: out = 32'b10000000000000000101110111100010; // input=-0.66943359375, output=-0.733446070462
			11'd1710: out = 32'b10000000000000000101111000001101; // input=-0.67041015625, output=-0.734761427651
			11'd1711: out = 32'b10000000000000000101111000111000; // input=-0.67138671875, output=-0.736078349955
			11'd1712: out = 32'b10000000000000000101111001100011; // input=-0.67236328125, output=-0.737396845268
			11'd1713: out = 32'b10000000000000000101111010001110; // input=-0.67333984375, output=-0.73871692154
			11'd1714: out = 32'b10000000000000000101111010111010; // input=-0.67431640625, output=-0.74003858678
			11'd1715: out = 32'b10000000000000000101111011100101; // input=-0.67529296875, output=-0.741361849058
			11'd1716: out = 32'b10000000000000000101111100010000; // input=-0.67626953125, output=-0.742686716502
			11'd1717: out = 32'b10000000000000000101111100111100; // input=-0.67724609375, output=-0.744013197301
			11'd1718: out = 32'b10000000000000000101111101100111; // input=-0.67822265625, output=-0.745341299708
			11'd1719: out = 32'b10000000000000000101111110010011; // input=-0.67919921875, output=-0.746671032034
			11'd1720: out = 32'b10000000000000000101111110111111; // input=-0.68017578125, output=-0.748002402655
			11'd1721: out = 32'b10000000000000000101111111101010; // input=-0.68115234375, output=-0.749335420011
			11'd1722: out = 32'b10000000000000000110000000010110; // input=-0.68212890625, output=-0.750670092604
			11'd1723: out = 32'b10000000000000000110000001000010; // input=-0.68310546875, output=-0.752006429003
			11'd1724: out = 32'b10000000000000000110000001101110; // input=-0.68408203125, output=-0.75334443784
			11'd1725: out = 32'b10000000000000000110000010011001; // input=-0.68505859375, output=-0.754684127815
			11'd1726: out = 32'b10000000000000000110000011000101; // input=-0.68603515625, output=-0.756025507694
			11'd1727: out = 32'b10000000000000000110000011110001; // input=-0.68701171875, output=-0.757368586311
			11'd1728: out = 32'b10000000000000000110000100011110; // input=-0.68798828125, output=-0.758713372569
			11'd1729: out = 32'b10000000000000000110000101001010; // input=-0.68896484375, output=-0.760059875439
			11'd1730: out = 32'b10000000000000000110000101110110; // input=-0.68994140625, output=-0.761408103962
			11'd1731: out = 32'b10000000000000000110000110100010; // input=-0.69091796875, output=-0.76275806725
			11'd1732: out = 32'b10000000000000000110000111001110; // input=-0.69189453125, output=-0.764109774486
			11'd1733: out = 32'b10000000000000000110000111111011; // input=-0.69287109375, output=-0.765463234926
			11'd1734: out = 32'b10000000000000000110001000100111; // input=-0.69384765625, output=-0.766818457899
			11'd1735: out = 32'b10000000000000000110001001010100; // input=-0.69482421875, output=-0.768175452807
			11'd1736: out = 32'b10000000000000000110001010000000; // input=-0.69580078125, output=-0.769534229128
			11'd1737: out = 32'b10000000000000000110001010101101; // input=-0.69677734375, output=-0.770894796414
			11'd1738: out = 32'b10000000000000000110001011011001; // input=-0.69775390625, output=-0.772257164294
			11'd1739: out = 32'b10000000000000000110001100000110; // input=-0.69873046875, output=-0.773621342475
			11'd1740: out = 32'b10000000000000000110001100110011; // input=-0.69970703125, output=-0.774987340742
			11'd1741: out = 32'b10000000000000000110001101100000; // input=-0.70068359375, output=-0.776355168958
			11'd1742: out = 32'b10000000000000000110001110001100; // input=-0.70166015625, output=-0.777724837066
			11'd1743: out = 32'b10000000000000000110001110111001; // input=-0.70263671875, output=-0.779096355093
			11'd1744: out = 32'b10000000000000000110001111100110; // input=-0.70361328125, output=-0.780469733143
			11'd1745: out = 32'b10000000000000000110010000010011; // input=-0.70458984375, output=-0.781844981407
			11'd1746: out = 32'b10000000000000000110010001000001; // input=-0.70556640625, output=-0.783222110157
			11'd1747: out = 32'b10000000000000000110010001101110; // input=-0.70654296875, output=-0.78460112975
			11'd1748: out = 32'b10000000000000000110010010011011; // input=-0.70751953125, output=-0.78598205063
			11'd1749: out = 32'b10000000000000000110010011001000; // input=-0.70849609375, output=-0.787364883328
			11'd1750: out = 32'b10000000000000000110010011110110; // input=-0.70947265625, output=-0.788749638461
			11'd1751: out = 32'b10000000000000000110010100100011; // input=-0.71044921875, output=-0.790136326735
			11'd1752: out = 32'b10000000000000000110010101010001; // input=-0.71142578125, output=-0.791524958947
			11'd1753: out = 32'b10000000000000000110010101111110; // input=-0.71240234375, output=-0.792915545985
			11'd1754: out = 32'b10000000000000000110010110101100; // input=-0.71337890625, output=-0.794308098827
			11'd1755: out = 32'b10000000000000000110010111011010; // input=-0.71435546875, output=-0.795702628547
			11'd1756: out = 32'b10000000000000000110011000000111; // input=-0.71533203125, output=-0.797099146312
			11'd1757: out = 32'b10000000000000000110011000110101; // input=-0.71630859375, output=-0.798497663382
			11'd1758: out = 32'b10000000000000000110011001100011; // input=-0.71728515625, output=-0.799898191117
			11'd1759: out = 32'b10000000000000000110011010010001; // input=-0.71826171875, output=-0.801300740973
			11'd1760: out = 32'b10000000000000000110011010111111; // input=-0.71923828125, output=-0.802705324505
			11'd1761: out = 32'b10000000000000000110011011101101; // input=-0.72021484375, output=-0.804111953369
			11'd1762: out = 32'b10000000000000000110011100011011; // input=-0.72119140625, output=-0.805520639322
			11'd1763: out = 32'b10000000000000000110011101001010; // input=-0.72216796875, output=-0.806931394221
			11'd1764: out = 32'b10000000000000000110011101111000; // input=-0.72314453125, output=-0.808344230032
			11'd1765: out = 32'b10000000000000000110011110100110; // input=-0.72412109375, output=-0.809759158821
			11'd1766: out = 32'b10000000000000000110011111010101; // input=-0.72509765625, output=-0.811176192763
			11'd1767: out = 32'b10000000000000000110100000000011; // input=-0.72607421875, output=-0.812595344141
			11'd1768: out = 32'b10000000000000000110100000110010; // input=-0.72705078125, output=-0.814016625347
			11'd1769: out = 32'b10000000000000000110100001100000; // input=-0.72802734375, output=-0.815440048882
			11'd1770: out = 32'b10000000000000000110100010001111; // input=-0.72900390625, output=-0.816865627361
			11'd1771: out = 32'b10000000000000000110100010111110; // input=-0.72998046875, output=-0.81829337351
			11'd1772: out = 32'b10000000000000000110100011101101; // input=-0.73095703125, output=-0.819723300173
			11'd1773: out = 32'b10000000000000000110100100011100; // input=-0.73193359375, output=-0.821155420307
			11'd1774: out = 32'b10000000000000000110100101001011; // input=-0.73291015625, output=-0.822589746989
			11'd1775: out = 32'b10000000000000000110100101111010; // input=-0.73388671875, output=-0.824026293413
			11'd1776: out = 32'b10000000000000000110100110101001; // input=-0.73486328125, output=-0.825465072897
			11'd1777: out = 32'b10000000000000000110100111011000; // input=-0.73583984375, output=-0.826906098877
			11'd1778: out = 32'b10000000000000000110101000000111; // input=-0.73681640625, output=-0.828349384918
			11'd1779: out = 32'b10000000000000000110101000110111; // input=-0.73779296875, output=-0.829794944707
			11'd1780: out = 32'b10000000000000000110101001100110; // input=-0.73876953125, output=-0.831242792059
			11'd1781: out = 32'b10000000000000000110101010010110; // input=-0.73974609375, output=-0.832692940918
			11'd1782: out = 32'b10000000000000000110101011000101; // input=-0.74072265625, output=-0.834145405359
			11'd1783: out = 32'b10000000000000000110101011110101; // input=-0.74169921875, output=-0.835600199588
			11'd1784: out = 32'b10000000000000000110101100100101; // input=-0.74267578125, output=-0.837057337948
			11'd1785: out = 32'b10000000000000000110101101010101; // input=-0.74365234375, output=-0.838516834915
			11'd1786: out = 32'b10000000000000000110101110000100; // input=-0.74462890625, output=-0.839978705103
			11'd1787: out = 32'b10000000000000000110101110110100; // input=-0.74560546875, output=-0.841442963267
			11'd1788: out = 32'b10000000000000000110101111100100; // input=-0.74658203125, output=-0.842909624303
			11'd1789: out = 32'b10000000000000000110110000010101; // input=-0.74755859375, output=-0.844378703249
			11'd1790: out = 32'b10000000000000000110110001000101; // input=-0.74853515625, output=-0.845850215289
			11'd1791: out = 32'b10000000000000000110110001110101; // input=-0.74951171875, output=-0.847324175756
			11'd1792: out = 32'b10000000000000000110110010100101; // input=-0.75048828125, output=-0.84880060013
			11'd1793: out = 32'b10000000000000000110110011010110; // input=-0.75146484375, output=-0.850279504044
			11'd1794: out = 32'b10000000000000000110110100000111; // input=-0.75244140625, output=-0.851760903282
			11'd1795: out = 32'b10000000000000000110110100110111; // input=-0.75341796875, output=-0.853244813787
			11'd1796: out = 32'b10000000000000000110110101101000; // input=-0.75439453125, output=-0.854731251657
			11'd1797: out = 32'b10000000000000000110110110011001; // input=-0.75537109375, output=-0.856220233152
			11'd1798: out = 32'b10000000000000000110110111001001; // input=-0.75634765625, output=-0.857711774692
			11'd1799: out = 32'b10000000000000000110110111111010; // input=-0.75732421875, output=-0.859205892863
			11'd1800: out = 32'b10000000000000000110111000101100; // input=-0.75830078125, output=-0.860702604419
			11'd1801: out = 32'b10000000000000000110111001011101; // input=-0.75927734375, output=-0.86220192628
			11'd1802: out = 32'b10000000000000000110111010001110; // input=-0.76025390625, output=-0.863703875539
			11'd1803: out = 32'b10000000000000000110111010111111; // input=-0.76123046875, output=-0.865208469465
			11'd1804: out = 32'b10000000000000000110111011110001; // input=-0.76220703125, output=-0.866715725501
			11'd1805: out = 32'b10000000000000000110111100100010; // input=-0.76318359375, output=-0.868225661271
			11'd1806: out = 32'b10000000000000000110111101010100; // input=-0.76416015625, output=-0.869738294579
			11'd1807: out = 32'b10000000000000000110111110000101; // input=-0.76513671875, output=-0.871253643414
			11'd1808: out = 32'b10000000000000000110111110110111; // input=-0.76611328125, output=-0.872771725953
			11'd1809: out = 32'b10000000000000000110111111101001; // input=-0.76708984375, output=-0.874292560562
			11'd1810: out = 32'b10000000000000000111000000011011; // input=-0.76806640625, output=-0.875816165799
			11'd1811: out = 32'b10000000000000000111000001001101; // input=-0.76904296875, output=-0.877342560418
			11'd1812: out = 32'b10000000000000000111000001111111; // input=-0.77001953125, output=-0.878871763373
			11'd1813: out = 32'b10000000000000000111000010110001; // input=-0.77099609375, output=-0.880403793817
			11'd1814: out = 32'b10000000000000000111000011100011; // input=-0.77197265625, output=-0.881938671108
			11'd1815: out = 32'b10000000000000000111000100010110; // input=-0.77294921875, output=-0.883476414811
			11'd1816: out = 32'b10000000000000000111000101001000; // input=-0.77392578125, output=-0.885017044704
			11'd1817: out = 32'b10000000000000000111000101111011; // input=-0.77490234375, output=-0.886560580776
			11'd1818: out = 32'b10000000000000000111000110101101; // input=-0.77587890625, output=-0.888107043235
			11'd1819: out = 32'b10000000000000000111000111100000; // input=-0.77685546875, output=-0.889656452506
			11'd1820: out = 32'b10000000000000000111001000010011; // input=-0.77783203125, output=-0.891208829243
			11'd1821: out = 32'b10000000000000000111001001000110; // input=-0.77880859375, output=-0.892764194322
			11'd1822: out = 32'b10000000000000000111001001111001; // input=-0.77978515625, output=-0.894322568854
			11'd1823: out = 32'b10000000000000000111001010101100; // input=-0.78076171875, output=-0.895883974181
			11'd1824: out = 32'b10000000000000000111001011100000; // input=-0.78173828125, output=-0.897448431885
			11'd1825: out = 32'b10000000000000000111001100010011; // input=-0.78271484375, output=-0.899015963789
			11'd1826: out = 32'b10000000000000000111001101000110; // input=-0.78369140625, output=-0.900586591962
			11'd1827: out = 32'b10000000000000000111001101111010; // input=-0.78466796875, output=-0.902160338722
			11'd1828: out = 32'b10000000000000000111001110101110; // input=-0.78564453125, output=-0.903737226641
			11'd1829: out = 32'b10000000000000000111001111100001; // input=-0.78662109375, output=-0.905317278548
			11'd1830: out = 32'b10000000000000000111010000010101; // input=-0.78759765625, output=-0.906900517533
			11'd1831: out = 32'b10000000000000000111010001001001; // input=-0.78857421875, output=-0.908486966953
			11'd1832: out = 32'b10000000000000000111010001111101; // input=-0.78955078125, output=-0.910076650436
			11'd1833: out = 32'b10000000000000000111010010110010; // input=-0.79052734375, output=-0.911669591883
			11'd1834: out = 32'b10000000000000000111010011100110; // input=-0.79150390625, output=-0.913265815473
			11'd1835: out = 32'b10000000000000000111010100011010; // input=-0.79248046875, output=-0.914865345673
			11'd1836: out = 32'b10000000000000000111010101001111; // input=-0.79345703125, output=-0.916468207233
			11'd1837: out = 32'b10000000000000000111010110000011; // input=-0.79443359375, output=-0.918074425201
			11'd1838: out = 32'b10000000000000000111010110111000; // input=-0.79541015625, output=-0.919684024919
			11'd1839: out = 32'b10000000000000000111010111101101; // input=-0.79638671875, output=-0.921297032036
			11'd1840: out = 32'b10000000000000000111011000100010; // input=-0.79736328125, output=-0.922913472506
			11'd1841: out = 32'b10000000000000000111011001010111; // input=-0.79833984375, output=-0.924533372597
			11'd1842: out = 32'b10000000000000000111011010001100; // input=-0.79931640625, output=-0.926156758898
			11'd1843: out = 32'b10000000000000000111011011000010; // input=-0.80029296875, output=-0.92778365832
			11'd1844: out = 32'b10000000000000000111011011110111; // input=-0.80126953125, output=-0.929414098105
			11'd1845: out = 32'b10000000000000000111011100101101; // input=-0.80224609375, output=-0.931048105828
			11'd1846: out = 32'b10000000000000000111011101100010; // input=-0.80322265625, output=-0.932685709409
			11'd1847: out = 32'b10000000000000000111011110011000; // input=-0.80419921875, output=-0.934326937112
			11'd1848: out = 32'b10000000000000000111011111001110; // input=-0.80517578125, output=-0.935971817557
			11'd1849: out = 32'b10000000000000000111100000000100; // input=-0.80615234375, output=-0.937620379721
			11'd1850: out = 32'b10000000000000000111100000111010; // input=-0.80712890625, output=-0.93927265295
			11'd1851: out = 32'b10000000000000000111100001110000; // input=-0.80810546875, output=-0.940928666959
			11'd1852: out = 32'b10000000000000000111100010100111; // input=-0.80908203125, output=-0.942588451845
			11'd1853: out = 32'b10000000000000000111100011011101; // input=-0.81005859375, output=-0.944252038088
			11'd1854: out = 32'b10000000000000000111100100010100; // input=-0.81103515625, output=-0.945919456565
			11'd1855: out = 32'b10000000000000000111100101001011; // input=-0.81201171875, output=-0.947590738548
			11'd1856: out = 32'b10000000000000000111100110000010; // input=-0.81298828125, output=-0.949265915721
			11'd1857: out = 32'b10000000000000000111100110111001; // input=-0.81396484375, output=-0.95094502018
			11'd1858: out = 32'b10000000000000000111100111110000; // input=-0.81494140625, output=-0.952628084445
			11'd1859: out = 32'b10000000000000000111101000100111; // input=-0.81591796875, output=-0.954315141464
			11'd1860: out = 32'b10000000000000000111101001011110; // input=-0.81689453125, output=-0.956006224626
			11'd1861: out = 32'b10000000000000000111101010010110; // input=-0.81787109375, output=-0.957701367765
			11'd1862: out = 32'b10000000000000000111101011001110; // input=-0.81884765625, output=-0.95940060517
			11'd1863: out = 32'b10000000000000000111101100000101; // input=-0.81982421875, output=-0.961103971595
			11'd1864: out = 32'b10000000000000000111101100111101; // input=-0.82080078125, output=-0.962811502264
			11'd1865: out = 32'b10000000000000000111101101110101; // input=-0.82177734375, output=-0.964523232885
			11'd1866: out = 32'b10000000000000000111101110101110; // input=-0.82275390625, output=-0.966239199654
			11'd1867: out = 32'b10000000000000000111101111100110; // input=-0.82373046875, output=-0.967959439271
			11'd1868: out = 32'b10000000000000000111110000011111; // input=-0.82470703125, output=-0.969683988941
			11'd1869: out = 32'b10000000000000000111110001010111; // input=-0.82568359375, output=-0.971412886393
			11'd1870: out = 32'b10000000000000000111110010010000; // input=-0.82666015625, output=-0.973146169884
			11'd1871: out = 32'b10000000000000000111110011001001; // input=-0.82763671875, output=-0.974883878213
			11'd1872: out = 32'b10000000000000000111110100000010; // input=-0.82861328125, output=-0.976626050731
			11'd1873: out = 32'b10000000000000000111110100111011; // input=-0.82958984375, output=-0.978372727348
			11'd1874: out = 32'b10000000000000000111110101110101; // input=-0.83056640625, output=-0.980123948551
			11'd1875: out = 32'b10000000000000000111110110101110; // input=-0.83154296875, output=-0.981879755413
			11'd1876: out = 32'b10000000000000000111110111101000; // input=-0.83251953125, output=-0.983640189601
			11'd1877: out = 32'b10000000000000000111111000100010; // input=-0.83349609375, output=-0.985405293394
			11'd1878: out = 32'b10000000000000000111111001011100; // input=-0.83447265625, output=-0.987175109694
			11'd1879: out = 32'b10000000000000000111111010010110; // input=-0.83544921875, output=-0.988949682035
			11'd1880: out = 32'b10000000000000000111111011010000; // input=-0.83642578125, output=-0.990729054601
			11'd1881: out = 32'b10000000000000000111111100001011; // input=-0.83740234375, output=-0.992513272239
			11'd1882: out = 32'b10000000000000000111111101000101; // input=-0.83837890625, output=-0.99430238047
			11'd1883: out = 32'b10000000000000000111111110000000; // input=-0.83935546875, output=-0.996096425507
			11'd1884: out = 32'b10000000000000000111111110111011; // input=-0.84033203125, output=-0.997895454266
			11'd1885: out = 32'b10000000000000000111111111110110; // input=-0.84130859375, output=-0.999699514384
			11'd1886: out = 32'b10000000000000001000000000110001; // input=-0.84228515625, output=-1.00150865423
			11'd1887: out = 32'b10000000000000001000000001101101; // input=-0.84326171875, output=-1.00332292294
			11'd1888: out = 32'b10000000000000001000000010101001; // input=-0.84423828125, output=-1.00514237039
			11'd1889: out = 32'b10000000000000001000000011100100; // input=-0.84521484375, output=-1.00696704727
			11'd1890: out = 32'b10000000000000001000000100100000; // input=-0.84619140625, output=-1.00879700506
			11'd1891: out = 32'b10000000000000001000000101011100; // input=-0.84716796875, output=-1.01063229605
			11'd1892: out = 32'b10000000000000001000000110011001; // input=-0.84814453125, output=-1.01247297339
			11'd1893: out = 32'b10000000000000001000000111010101; // input=-0.84912109375, output=-1.01431909107
			11'd1894: out = 32'b10000000000000001000001000010010; // input=-0.85009765625, output=-1.01617070397
			11'd1895: out = 32'b10000000000000001000001001001111; // input=-0.85107421875, output=-1.01802786786
			11'd1896: out = 32'b10000000000000001000001010001100; // input=-0.85205078125, output=-1.01989063942
			11'd1897: out = 32'b10000000000000001000001011001001; // input=-0.85302734375, output=-1.02175907629
			11'd1898: out = 32'b10000000000000001000001100000110; // input=-0.85400390625, output=-1.02363323705
			11'd1899: out = 32'b10000000000000001000001101000100; // input=-0.85498046875, output=-1.02551318129
			11'd1900: out = 32'b10000000000000001000001110000010; // input=-0.85595703125, output=-1.02739896957
			11'd1901: out = 32'b10000000000000001000001111000000; // input=-0.85693359375, output=-1.02929066351
			11'd1902: out = 32'b10000000000000001000001111111110; // input=-0.85791015625, output=-1.03118832579
			11'd1903: out = 32'b10000000000000001000010000111100; // input=-0.85888671875, output=-1.03309202014
			11'd1904: out = 32'b10000000000000001000010001111011; // input=-0.85986328125, output=-1.03500181142
			11'd1905: out = 32'b10000000000000001000010010111010; // input=-0.86083984375, output=-1.03691776563
			11'd1906: out = 32'b10000000000000001000010011111001; // input=-0.86181640625, output=-1.03883994992
			11'd1907: out = 32'b10000000000000001000010100111000; // input=-0.86279296875, output=-1.04076843263
			11'd1908: out = 32'b10000000000000001000010101110111; // input=-0.86376953125, output=-1.04270328333
			11'd1909: out = 32'b10000000000000001000010110110111; // input=-0.86474609375, output=-1.04464457284
			11'd1910: out = 32'b10000000000000001000010111110111; // input=-0.86572265625, output=-1.04659237326
			11'd1911: out = 32'b10000000000000001000011000110111; // input=-0.86669921875, output=-1.04854675801
			11'd1912: out = 32'b10000000000000001000011001110111; // input=-0.86767578125, output=-1.05050780186
			11'd1913: out = 32'b10000000000000001000011010111000; // input=-0.86865234375, output=-1.05247558096
			11'd1914: out = 32'b10000000000000001000011011111000; // input=-0.86962890625, output=-1.0544501729
			11'd1915: out = 32'b10000000000000001000011100111001; // input=-0.87060546875, output=-1.0564316567
			11'd1916: out = 32'b10000000000000001000011101111010; // input=-0.87158203125, output=-1.0584201129
			11'd1917: out = 32'b10000000000000001000011110111100; // input=-0.87255859375, output=-1.06041562356
			11'd1918: out = 32'b10000000000000001000011111111101; // input=-0.87353515625, output=-1.06241827236
			11'd1919: out = 32'b10000000000000001000100000111111; // input=-0.87451171875, output=-1.06442814454
			11'd1920: out = 32'b10000000000000001000100010000001; // input=-0.87548828125, output=-1.06644532706
			11'd1921: out = 32'b10000000000000001000100011000100; // input=-0.87646484375, output=-1.06846990857
			11'd1922: out = 32'b10000000000000001000100100000110; // input=-0.87744140625, output=-1.07050197947
			11'd1923: out = 32'b10000000000000001000100101001001; // input=-0.87841796875, output=-1.07254163199
			11'd1924: out = 32'b10000000000000001000100110001100; // input=-0.87939453125, output=-1.0745889602
			11'd1925: out = 32'b10000000000000001000100111001111; // input=-0.88037109375, output=-1.07664406011
			11'd1926: out = 32'b10000000000000001000101000010011; // input=-0.88134765625, output=-1.07870702967
			11'd1927: out = 32'b10000000000000001000101001010111; // input=-0.88232421875, output=-1.08077796888
			11'd1928: out = 32'b10000000000000001000101010011011; // input=-0.88330078125, output=-1.08285697979
			11'd1929: out = 32'b10000000000000001000101011011111; // input=-0.88427734375, output=-1.08494416663
			11'd1930: out = 32'b10000000000000001000101100100100; // input=-0.88525390625, output=-1.08703963583
			11'd1931: out = 32'b10000000000000001000101101101001; // input=-0.88623046875, output=-1.08914349607
			11'd1932: out = 32'b10000000000000001000101110101110; // input=-0.88720703125, output=-1.09125585841
			11'd1933: out = 32'b10000000000000001000101111110100; // input=-0.88818359375, output=-1.09337683631
			11'd1934: out = 32'b10000000000000001000110000111010; // input=-0.88916015625, output=-1.0955065457
			11'd1935: out = 32'b10000000000000001000110010000000; // input=-0.89013671875, output=-1.0976451051
			11'd1936: out = 32'b10000000000000001000110011000110; // input=-0.89111328125, output=-1.09979263568
			11'd1937: out = 32'b10000000000000001000110100001101; // input=-0.89208984375, output=-1.10194926132
			11'd1938: out = 32'b10000000000000001000110101010100; // input=-0.89306640625, output=-1.10411510871
			11'd1939: out = 32'b10000000000000001000110110011011; // input=-0.89404296875, output=-1.10629030749
			11'd1940: out = 32'b10000000000000001000110111100011; // input=-0.89501953125, output=-1.10847499025
			11'd1941: out = 32'b10000000000000001000111000101010; // input=-0.89599609375, output=-1.1106692927
			11'd1942: out = 32'b10000000000000001000111001110011; // input=-0.89697265625, output=-1.11287335376
			11'd1943: out = 32'b10000000000000001000111010111011; // input=-0.89794921875, output=-1.11508731565
			11'd1944: out = 32'b10000000000000001000111100000100; // input=-0.89892578125, output=-1.117311324
			11'd1945: out = 32'b10000000000000001000111101001101; // input=-0.89990234375, output=-1.11954552799
			11'd1946: out = 32'b10000000000000001000111110010111; // input=-0.90087890625, output=-1.12179008044
			11'd1947: out = 32'b10000000000000001000111111100001; // input=-0.90185546875, output=-1.12404513797
			11'd1948: out = 32'b10000000000000001001000000101011; // input=-0.90283203125, output=-1.1263108611
			11'd1949: out = 32'b10000000000000001001000001110110; // input=-0.90380859375, output=-1.12858741441
			11'd1950: out = 32'b10000000000000001001000011000001; // input=-0.90478515625, output=-1.13087496667
			11'd1951: out = 32'b10000000000000001001000100001100; // input=-0.90576171875, output=-1.13317369102
			11'd1952: out = 32'b10000000000000001001000101011000; // input=-0.90673828125, output=-1.13548376509
			11'd1953: out = 32'b10000000000000001001000110100100; // input=-0.90771484375, output=-1.13780537118
			11'd1954: out = 32'b10000000000000001001000111110000; // input=-0.90869140625, output=-1.14013869645
			11'd1955: out = 32'b10000000000000001001001000111101; // input=-0.90966796875, output=-1.14248393307
			11'd1956: out = 32'b10000000000000001001001010001010; // input=-0.91064453125, output=-1.14484127846
			11'd1957: out = 32'b10000000000000001001001011011000; // input=-0.91162109375, output=-1.14721093543
			11'd1958: out = 32'b10000000000000001001001100100110; // input=-0.91259765625, output=-1.14959311244
			11'd1959: out = 32'b10000000000000001001001101110100; // input=-0.91357421875, output=-1.1519880238
			11'd1960: out = 32'b10000000000000001001001111000011; // input=-0.91455078125, output=-1.1543958899
			11'd1961: out = 32'b10000000000000001001010000010011; // input=-0.91552734375, output=-1.15681693745
			11'd1962: out = 32'b10000000000000001001010001100010; // input=-0.91650390625, output=-1.15925139978
			11'd1963: out = 32'b10000000000000001001010010110011; // input=-0.91748046875, output=-1.16169951703
			11'd1964: out = 32'b10000000000000001001010100000011; // input=-0.91845703125, output=-1.16416153653
			11'd1965: out = 32'b10000000000000001001010101010100; // input=-0.91943359375, output=-1.16663771301
			11'd1966: out = 32'b10000000000000001001010110100110; // input=-0.92041015625, output=-1.16912830899
			11'd1967: out = 32'b10000000000000001001010111111000; // input=-0.92138671875, output=-1.17163359507
			11'd1968: out = 32'b10000000000000001001011001001011; // input=-0.92236328125, output=-1.17415385031
			11'd1969: out = 32'b10000000000000001001011010011110; // input=-0.92333984375, output=-1.17668936258
			11'd1970: out = 32'b10000000000000001001011011110001; // input=-0.92431640625, output=-1.17924042897
			11'd1971: out = 32'b10000000000000001001011101000101; // input=-0.92529296875, output=-1.18180735621
			11'd1972: out = 32'b10000000000000001001011110011010; // input=-0.92626953125, output=-1.1843904611
			11'd1973: out = 32'b10000000000000001001011111101111; // input=-0.92724609375, output=-1.18699007099
			11'd1974: out = 32'b10000000000000001001100001000101; // input=-0.92822265625, output=-1.18960652428
			11'd1975: out = 32'b10000000000000001001100010011011; // input=-0.92919921875, output=-1.19224017094
			11'd1976: out = 32'b10000000000000001001100011110010; // input=-0.93017578125, output=-1.19489137306
			11'd1977: out = 32'b10000000000000001001100101001010; // input=-0.93115234375, output=-1.1975605055
			11'd1978: out = 32'b10000000000000001001100110100010; // input=-0.93212890625, output=-1.20024795643
			11'd1979: out = 32'b10000000000000001001100111111010; // input=-0.93310546875, output=-1.20295412811
			11'd1980: out = 32'b10000000000000001001101001010100; // input=-0.93408203125, output=-1.20567943755
			11'd1981: out = 32'b10000000000000001001101010101110; // input=-0.93505859375, output=-1.20842431728
			11'd1982: out = 32'b10000000000000001001101100001000; // input=-0.93603515625, output=-1.21118921619
			11'd1983: out = 32'b10000000000000001001101101100100; // input=-0.93701171875, output=-1.2139746004
			11'd1984: out = 32'b10000000000000001001101110111111; // input=-0.93798828125, output=-1.21678095422
			11'd1985: out = 32'b10000000000000001001110000011100; // input=-0.93896484375, output=-1.21960878111
			11'd1986: out = 32'b10000000000000001001110001111010; // input=-0.93994140625, output=-1.22245860481
			11'd1987: out = 32'b10000000000000001001110011011000; // input=-0.94091796875, output=-1.22533097047
			11'd1988: out = 32'b10000000000000001001110100110111; // input=-0.94189453125, output=-1.22822644589
			11'd1989: out = 32'b10000000000000001001110110010110; // input=-0.94287109375, output=-1.23114562288
			11'd1990: out = 32'b10000000000000001001110111110111; // input=-0.94384765625, output=-1.23408911871
			11'd1991: out = 32'b10000000000000001001111001011000; // input=-0.94482421875, output=-1.23705757763
			11'd1992: out = 32'b10000000000000001001111010111010; // input=-0.94580078125, output=-1.24005167258
			11'd1993: out = 32'b10000000000000001001111100011101; // input=-0.94677734375, output=-1.24307210702
			11'd1994: out = 32'b10000000000000001001111110000001; // input=-0.94775390625, output=-1.24611961686
			11'd1995: out = 32'b10000000000000001001111111100110; // input=-0.94873046875, output=-1.24919497264
			11'd1996: out = 32'b10000000000000001010000001001011; // input=-0.94970703125, output=-1.25229898181
			11'd1997: out = 32'b10000000000000001010000010110010; // input=-0.95068359375, output=-1.25543249128
			11'd1998: out = 32'b10000000000000001010000100011010; // input=-0.95166015625, output=-1.25859639018
			11'd1999: out = 32'b10000000000000001010000110000010; // input=-0.95263671875, output=-1.26179161284
			11'd2000: out = 32'b10000000000000001010000111101100; // input=-0.95361328125, output=-1.26501914206
			11'd2001: out = 32'b10000000000000001010001001010111; // input=-0.95458984375, output=-1.26828001276
			11'd2002: out = 32'b10000000000000001010001011000011; // input=-0.95556640625, output=-1.27157531586
			11'd2003: out = 32'b10000000000000001010001100110000; // input=-0.95654296875, output=-1.27490620266
			11'd2004: out = 32'b10000000000000001010001110011110; // input=-0.95751953125, output=-1.27827388961
			11'd2005: out = 32'b10000000000000001010010000001110; // input=-0.95849609375, output=-1.28167966359
			11'd2006: out = 32'b10000000000000001010010001111111; // input=-0.95947265625, output=-1.28512488772
			11'd2007: out = 32'b10000000000000001010010011110001; // input=-0.96044921875, output=-1.28861100788
			11'd2008: out = 32'b10000000000000001010010101100101; // input=-0.96142578125, output=-1.2921395599
			11'd2009: out = 32'b10000000000000001010010111011010; // input=-0.96240234375, output=-1.29571217755
			11'd2010: out = 32'b10000000000000001010011001010000; // input=-0.96337890625, output=-1.29933060156
			11'd2011: out = 32'b10000000000000001010011011001001; // input=-0.96435546875, output=-1.30299668967
			11'd2012: out = 32'b10000000000000001010011101000010; // input=-0.96533203125, output=-1.30671242792
			11'd2013: out = 32'b10000000000000001010011110111110; // input=-0.96630859375, output=-1.3104799434
			11'd2014: out = 32'b10000000000000001010100000111011; // input=-0.96728515625, output=-1.31430151869
			11'd2015: out = 32'b10000000000000001010100010111010; // input=-0.96826171875, output=-1.31817960826
			11'd2016: out = 32'b10000000000000001010100100111011; // input=-0.96923828125, output=-1.32211685711
			11'd2017: out = 32'b10000000000000001010100110111110; // input=-0.97021484375, output=-1.32611612215
			11'd2018: out = 32'b10000000000000001010101001000011; // input=-0.97119140625, output=-1.33018049673
			11'd2019: out = 32'b10000000000000001010101011001011; // input=-0.97216796875, output=-1.33431333899
			11'd2020: out = 32'b10000000000000001010101101010101; // input=-0.97314453125, output=-1.33851830468
			11'd2021: out = 32'b10000000000000001010101111100001; // input=-0.97412109375, output=-1.34279938541
			11'd2022: out = 32'b10000000000000001010110001110000; // input=-0.97509765625, output=-1.34716095354
			11'd2023: out = 32'b10000000000000001010110100000001; // input=-0.97607421875, output=-1.35160781497
			11'd2024: out = 32'b10000000000000001010110110010110; // input=-0.97705078125, output=-1.35614527182
			11'd2025: out = 32'b10000000000000001010111000101110; // input=-0.97802734375, output=-1.36077919721
			11'd2026: out = 32'b10000000000000001010111011001001; // input=-0.97900390625, output=-1.36551612523
			11'd2027: out = 32'b10000000000000001010111101101000; // input=-0.97998046875, output=-1.37036335996
			11'd2028: out = 32'b10000000000000001011000000001011; // input=-0.98095703125, output=-1.37532910873
			11'd2029: out = 32'b10000000000000001011000010110010; // input=-0.98193359375, output=-1.38042264672
			11'd2030: out = 32'b10000000000000001011000101011101; // input=-0.98291015625, output=-1.38565452202
			11'd2031: out = 32'b10000000000000001011001000001101; // input=-0.98388671875, output=-1.39103681451
			11'd2032: out = 32'b10000000000000001011001011000011; // input=-0.98486328125, output=-1.39658346647
			11'd2033: out = 32'b10000000000000001011001101111111; // input=-0.98583984375, output=-1.40231071107
			11'd2034: out = 32'b10000000000000001011010001000001; // input=-0.98681640625, output=-1.40823763659
			11'd2035: out = 32'b10000000000000001011010100001011; // input=-0.98779296875, output=-1.41438694293
			11'd2036: out = 32'b10000000000000001011010111011100; // input=-0.98876953125, output=-1.42078597714
			11'd2037: out = 32'b10000000000000001011011010110111; // input=-0.98974609375, output=-1.42746818517
			11'd2038: out = 32'b10000000000000001011011110011101; // input=-0.99072265625, output=-1.43447520447
			11'd2039: out = 32'b10000000000000001011100010001111; // input=-0.99169921875, output=-1.44185998152
			11'd2040: out = 32'b10000000000000001011100110001111; // input=-0.99267578125, output=-1.44969160393
			11'd2041: out = 32'b10000000000000001011101010100010; // input=-0.99365234375, output=-1.45806316311
			11'd2042: out = 32'b10000000000000001011101111001010; // input=-0.99462890625, output=-1.46710535557
			11'd2043: out = 32'b10000000000000001011110100001111; // input=-0.99560546875, output=-1.47701196053
			11'd2044: out = 32'b10000000000000001011111001111010; // input=-0.99658203125, output=-1.48809303047
			11'd2045: out = 32'b10000000000000001100000000011110; // input=-0.99755859375, output=-1.50090497815
			11'd2046: out = 32'b10000000000000001100001000100010; // input=-0.99853515625, output=-1.51666312963
			11'd2047: out = 32'b10000000000000001100010100010000; // input=-0.99951171875, output=-1.53954505509
		endcase
	end
	converter_arc U0 (a, index);

endmodule

module converter_arc(a, index);
	input  [31:0] a;
	output [10:0] index;
	assign index[10]   = a[31];
	assign index[9:0]  = (a[15]) ? 10'b1111111111 : a[14:5];
endmodule
