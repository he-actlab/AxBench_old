// Developed by: Amir Yazdanbakhsh
// Email: a.yazdanbakhsh@gatech.edu

`timescale 1ns/1ps
module cos_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000000111111111111111; // input=0.001953125, output=0.999998092652
			11'd1: out = 32'b00000000000000000111111111111111; // input=0.005859375, output=0.999982833911
			11'd2: out = 32'b00000000000000000111111111111110; // input=0.009765625, output=0.999952316663
			11'd3: out = 32'b00000000000000000111111111111101; // input=0.013671875, output=0.999906541373
			11'd4: out = 32'b00000000000000000111111111111011; // input=0.017578125, output=0.999845508739
			11'd5: out = 32'b00000000000000000111111111111000; // input=0.021484375, output=0.999769219693
			11'd6: out = 32'b00000000000000000111111111110101; // input=0.025390625, output=0.999677675398
			11'd7: out = 32'b00000000000000000111111111110010; // input=0.029296875, output=0.999570877252
			11'd8: out = 32'b00000000000000000111111111101110; // input=0.033203125, output=0.999448826885
			11'd9: out = 32'b00000000000000000111111111101001; // input=0.037109375, output=0.999311526157
			11'd10: out = 32'b00000000000000000111111111100100; // input=0.041015625, output=0.999158977166
			11'd11: out = 32'b00000000000000000111111111011111; // input=0.044921875, output=0.998991182238
			11'd12: out = 32'b00000000000000000111111111011001; // input=0.048828125, output=0.998808143933
			11'd13: out = 32'b00000000000000000111111111010010; // input=0.052734375, output=0.998609865045
			11'd14: out = 32'b00000000000000000111111111001011; // input=0.056640625, output=0.998396348599
			11'd15: out = 32'b00000000000000000111111111000100; // input=0.060546875, output=0.998167597854
			11'd16: out = 32'b00000000000000000111111110111100; // input=0.064453125, output=0.997923616299
			11'd17: out = 32'b00000000000000000111111110110011; // input=0.068359375, output=0.997664407657
			11'd18: out = 32'b00000000000000000111111110101010; // input=0.072265625, output=0.997389975884
			11'd19: out = 32'b00000000000000000111111110100001; // input=0.076171875, output=0.997100325166
			11'd20: out = 32'b00000000000000000111111110010111; // input=0.080078125, output=0.996795459925
			11'd21: out = 32'b00000000000000000111111110001101; // input=0.083984375, output=0.996475384812
			11'd22: out = 32'b00000000000000000111111110000010; // input=0.087890625, output=0.99614010471
			11'd23: out = 32'b00000000000000000111111101110110; // input=0.091796875, output=0.995789624735
			11'd24: out = 32'b00000000000000000111111101101010; // input=0.095703125, output=0.995423950236
			11'd25: out = 32'b00000000000000000111111101011110; // input=0.099609375, output=0.995043086793
			11'd26: out = 32'b00000000000000000111111101010001; // input=0.103515625, output=0.994647040216
			11'd27: out = 32'b00000000000000000111111101000011; // input=0.107421875, output=0.994235816549
			11'd28: out = 32'b00000000000000000111111100110101; // input=0.111328125, output=0.993809422066
			11'd29: out = 32'b00000000000000000111111100100111; // input=0.115234375, output=0.993367863275
			11'd30: out = 32'b00000000000000000111111100011000; // input=0.119140625, output=0.992911146912
			11'd31: out = 32'b00000000000000000111111100001000; // input=0.123046875, output=0.992439279947
			11'd32: out = 32'b00000000000000000111111011111000; // input=0.126953125, output=0.991952269579
			11'd33: out = 32'b00000000000000000111111011101000; // input=0.130859375, output=0.99145012324
			11'd34: out = 32'b00000000000000000111111011010111; // input=0.134765625, output=0.990932848592
			11'd35: out = 32'b00000000000000000111111011000101; // input=0.138671875, output=0.990400453528
			11'd36: out = 32'b00000000000000000111111010110100; // input=0.142578125, output=0.989852946172
			11'd37: out = 32'b00000000000000000111111010100001; // input=0.146484375, output=0.989290334878
			11'd38: out = 32'b00000000000000000111111010001110; // input=0.150390625, output=0.98871262823
			11'd39: out = 32'b00000000000000000111111001111011; // input=0.154296875, output=0.988119835044
			11'd40: out = 32'b00000000000000000111111001100111; // input=0.158203125, output=0.987511964365
			11'd41: out = 32'b00000000000000000111111001010010; // input=0.162109375, output=0.986889025468
			11'd42: out = 32'b00000000000000000111111000111101; // input=0.166015625, output=0.986251027859
			11'd43: out = 32'b00000000000000000111111000101000; // input=0.169921875, output=0.985597981273
			11'd44: out = 32'b00000000000000000111111000010010; // input=0.173828125, output=0.984929895674
			11'd45: out = 32'b00000000000000000111110111111100; // input=0.177734375, output=0.984246781257
			11'd46: out = 32'b00000000000000000111110111100101; // input=0.181640625, output=0.983548648445
			11'd47: out = 32'b00000000000000000111110111001110; // input=0.185546875, output=0.98283550789
			11'd48: out = 32'b00000000000000000111110110110110; // input=0.189453125, output=0.982107370475
			11'd49: out = 32'b00000000000000000111110110011101; // input=0.193359375, output=0.98136424731
			11'd50: out = 32'b00000000000000000111110110000101; // input=0.197265625, output=0.980606149734
			11'd51: out = 32'b00000000000000000111110101101011; // input=0.201171875, output=0.979833089314
			11'd52: out = 32'b00000000000000000111110101010001; // input=0.205078125, output=0.979045077847
			11'd53: out = 32'b00000000000000000111110100110111; // input=0.208984375, output=0.978242127357
			11'd54: out = 32'b00000000000000000111110100011100; // input=0.212890625, output=0.977424250095
			11'd55: out = 32'b00000000000000000111110100000001; // input=0.216796875, output=0.976591458542
			11'd56: out = 32'b00000000000000000111110011100101; // input=0.220703125, output=0.975743765405
			11'd57: out = 32'b00000000000000000111110011001001; // input=0.224609375, output=0.974881183619
			11'd58: out = 32'b00000000000000000111110010101100; // input=0.228515625, output=0.974003726345
			11'd59: out = 32'b00000000000000000111110010001111; // input=0.232421875, output=0.973111406972
			11'd60: out = 32'b00000000000000000111110001110001; // input=0.236328125, output=0.972204239117
			11'd61: out = 32'b00000000000000000111110001010011; // input=0.240234375, output=0.971282236621
			11'd62: out = 32'b00000000000000000111110000110100; // input=0.244140625, output=0.970345413553
			11'd63: out = 32'b00000000000000000111110000010101; // input=0.248046875, output=0.969393784208
			11'd64: out = 32'b00000000000000000111101111110101; // input=0.251953125, output=0.968427363107
			11'd65: out = 32'b00000000000000000111101111010101; // input=0.255859375, output=0.967446164995
			11'd66: out = 32'b00000000000000000111101110110101; // input=0.259765625, output=0.966450204846
			11'd67: out = 32'b00000000000000000111101110010100; // input=0.263671875, output=0.965439497855
			11'd68: out = 32'b00000000000000000111101101110010; // input=0.267578125, output=0.964414059445
			11'd69: out = 32'b00000000000000000111101101010000; // input=0.271484375, output=0.963373905264
			11'd70: out = 32'b00000000000000000111101100101101; // input=0.275390625, output=0.962319051181
			11'd71: out = 32'b00000000000000000111101100001010; // input=0.279296875, output=0.961249513295
			11'd72: out = 32'b00000000000000000111101011100111; // input=0.283203125, output=0.960165307923
			11'd73: out = 32'b00000000000000000111101011000011; // input=0.287109375, output=0.95906645161
			11'd74: out = 32'b00000000000000000111101010011110; // input=0.291015625, output=0.957952961123
			11'd75: out = 32'b00000000000000000111101001111001; // input=0.294921875, output=0.956824853452
			11'd76: out = 32'b00000000000000000111101001010100; // input=0.298828125, output=0.955682145811
			11'd77: out = 32'b00000000000000000111101000101110; // input=0.302734375, output=0.954524855637
			11'd78: out = 32'b00000000000000000111101000000111; // input=0.306640625, output=0.953353000587
			11'd79: out = 32'b00000000000000000111100111100001; // input=0.310546875, output=0.952166598544
			11'd80: out = 32'b00000000000000000111100110111001; // input=0.314453125, output=0.95096566761
			11'd81: out = 32'b00000000000000000111100110010001; // input=0.318359375, output=0.94975022611
			11'd82: out = 32'b00000000000000000111100101101001; // input=0.322265625, output=0.94852029259
			11'd83: out = 32'b00000000000000000111100101000000; // input=0.326171875, output=0.947275885817
			11'd84: out = 32'b00000000000000000111100100010111; // input=0.330078125, output=0.94601702478
			11'd85: out = 32'b00000000000000000111100011101101; // input=0.333984375, output=0.944743728687
			11'd86: out = 32'b00000000000000000111100011000011; // input=0.337890625, output=0.943456016966
			11'd87: out = 32'b00000000000000000111100010011000; // input=0.341796875, output=0.942153909268
			11'd88: out = 32'b00000000000000000111100001101101; // input=0.345703125, output=0.940837425461
			11'd89: out = 32'b00000000000000000111100001000010; // input=0.349609375, output=0.939506585632
			11'd90: out = 32'b00000000000000000111100000010110; // input=0.353515625, output=0.938161410088
			11'd91: out = 32'b00000000000000000111011111101001; // input=0.357421875, output=0.936801919355
			11'd92: out = 32'b00000000000000000111011110111100; // input=0.361328125, output=0.935428134178
			11'd93: out = 32'b00000000000000000111011110001111; // input=0.365234375, output=0.934040075518
			11'd94: out = 32'b00000000000000000111011101100001; // input=0.369140625, output=0.932637764556
			11'd95: out = 32'b00000000000000000111011100110010; // input=0.373046875, output=0.931221222689
			11'd96: out = 32'b00000000000000000111011100000011; // input=0.376953125, output=0.929790471532
			11'd97: out = 32'b00000000000000000111011011010100; // input=0.380859375, output=0.928345532916
			11'd98: out = 32'b00000000000000000111011010100100; // input=0.384765625, output=0.92688642889
			11'd99: out = 32'b00000000000000000111011001110100; // input=0.388671875, output=0.925413181717
			11'd100: out = 32'b00000000000000000111011001000011; // input=0.392578125, output=0.923925813877
			11'd101: out = 32'b00000000000000000111011000010010; // input=0.396484375, output=0.922424348067
			11'd102: out = 32'b00000000000000000111010111100000; // input=0.400390625, output=0.920908807195
			11'd103: out = 32'b00000000000000000111010110101110; // input=0.404296875, output=0.919379214389
			11'd104: out = 32'b00000000000000000111010101111100; // input=0.408203125, output=0.917835592986
			11'd105: out = 32'b00000000000000000111010101001001; // input=0.412109375, output=0.916277966542
			11'd106: out = 32'b00000000000000000111010100010101; // input=0.416015625, output=0.914706358823
			11'd107: out = 32'b00000000000000000111010011100001; // input=0.419921875, output=0.913120793811
			11'd108: out = 32'b00000000000000000111010010101101; // input=0.423828125, output=0.911521295699
			11'd109: out = 32'b00000000000000000111010001111000; // input=0.427734375, output=0.909907888893
			11'd110: out = 32'b00000000000000000111010001000011; // input=0.431640625, output=0.908280598013
			11'd111: out = 32'b00000000000000000111010000001101; // input=0.435546875, output=0.906639447888
			11'd112: out = 32'b00000000000000000111001111010111; // input=0.439453125, output=0.90498446356
			11'd113: out = 32'b00000000000000000111001110100000; // input=0.443359375, output=0.903315670283
			11'd114: out = 32'b00000000000000000111001101101001; // input=0.447265625, output=0.901633093521
			11'd115: out = 32'b00000000000000000111001100110001; // input=0.451171875, output=0.899936758946
			11'd116: out = 32'b00000000000000000111001011111001; // input=0.455078125, output=0.898226692444
			11'd117: out = 32'b00000000000000000111001011000001; // input=0.458984375, output=0.896502920108
			11'd118: out = 32'b00000000000000000111001010001000; // input=0.462890625, output=0.89476546824
			11'd119: out = 32'b00000000000000000111001001001110; // input=0.466796875, output=0.893014363352
			11'd120: out = 32'b00000000000000000111001000010100; // input=0.470703125, output=0.891249632163
			11'd121: out = 32'b00000000000000000111000111011010; // input=0.474609375, output=0.889471301602
			11'd122: out = 32'b00000000000000000111000110011111; // input=0.478515625, output=0.887679398803
			11'd123: out = 32'b00000000000000000111000101100100; // input=0.482421875, output=0.885873951108
			11'd124: out = 32'b00000000000000000111000100101001; // input=0.486328125, output=0.884054986067
			11'd125: out = 32'b00000000000000000111000011101101; // input=0.490234375, output=0.882222531435
			11'd126: out = 32'b00000000000000000111000010110000; // input=0.494140625, output=0.880376615172
			11'd127: out = 32'b00000000000000000111000001110011; // input=0.498046875, output=0.878517265445
			11'd128: out = 32'b00000000000000000111000000110110; // input=0.501953125, output=0.876644510625
			11'd129: out = 32'b00000000000000000110111111111000; // input=0.505859375, output=0.874758379289
			11'd130: out = 32'b00000000000000000110111110111010; // input=0.509765625, output=0.872858900216
			11'd131: out = 32'b00000000000000000110111101111011; // input=0.513671875, output=0.870946102391
			11'd132: out = 32'b00000000000000000110111100111100; // input=0.517578125, output=0.869020014999
			11'd133: out = 32'b00000000000000000110111011111100; // input=0.521484375, output=0.867080667431
			11'd134: out = 32'b00000000000000000110111010111101; // input=0.525390625, output=0.865128089279
			11'd135: out = 32'b00000000000000000110111001111100; // input=0.529296875, output=0.863162310337
			11'd136: out = 32'b00000000000000000110111000111011; // input=0.533203125, output=0.861183360599
			11'd137: out = 32'b00000000000000000110110111111010; // input=0.537109375, output=0.859191270264
			11'd138: out = 32'b00000000000000000110110110111000; // input=0.541015625, output=0.857186069726
			11'd139: out = 32'b00000000000000000110110101110110; // input=0.544921875, output=0.855167789584
			11'd140: out = 32'b00000000000000000110110100110100; // input=0.548828125, output=0.853136460634
			11'd141: out = 32'b00000000000000000110110011110001; // input=0.552734375, output=0.85109211387
			11'd142: out = 32'b00000000000000000110110010101101; // input=0.556640625, output=0.849034780489
			11'd143: out = 32'b00000000000000000110110001101001; // input=0.560546875, output=0.846964491881
			11'd144: out = 32'b00000000000000000110110000100101; // input=0.564453125, output=0.844881279637
			11'd145: out = 32'b00000000000000000110101111100000; // input=0.568359375, output=0.842785175544
			11'd146: out = 32'b00000000000000000110101110011011; // input=0.572265625, output=0.840676211586
			11'd147: out = 32'b00000000000000000110101101010110; // input=0.576171875, output=0.838554419944
			11'd148: out = 32'b00000000000000000110101100010000; // input=0.580078125, output=0.836419832992
			11'd149: out = 32'b00000000000000000110101011001001; // input=0.583984375, output=0.834272483304
			11'd150: out = 32'b00000000000000000110101010000011; // input=0.587890625, output=0.832112403643
			11'd151: out = 32'b00000000000000000110101000111011; // input=0.591796875, output=0.829939626972
			11'd152: out = 32'b00000000000000000110100111110100; // input=0.595703125, output=0.827754186442
			11'd153: out = 32'b00000000000000000110100110101100; // input=0.599609375, output=0.825556115402
			11'd154: out = 32'b00000000000000000110100101100011; // input=0.603515625, output=0.823345447392
			11'd155: out = 32'b00000000000000000110100100011011; // input=0.607421875, output=0.821122216143
			11'd156: out = 32'b00000000000000000110100011010001; // input=0.611328125, output=0.818886455579
			11'd157: out = 32'b00000000000000000110100010001000; // input=0.615234375, output=0.816638199815
			11'd158: out = 32'b00000000000000000110100000111110; // input=0.619140625, output=0.814377483157
			11'd159: out = 32'b00000000000000000110011111110011; // input=0.623046875, output=0.812104340101
			11'd160: out = 32'b00000000000000000110011110101000; // input=0.626953125, output=0.809818805332
			11'd161: out = 32'b00000000000000000110011101011101; // input=0.630859375, output=0.807520913724
			11'd162: out = 32'b00000000000000000110011100010001; // input=0.634765625, output=0.80521070034
			11'd163: out = 32'b00000000000000000110011011000101; // input=0.638671875, output=0.802888200432
			11'd164: out = 32'b00000000000000000110011001111001; // input=0.642578125, output=0.800553449438
			11'd165: out = 32'b00000000000000000110011000101100; // input=0.646484375, output=0.798206482983
			11'd166: out = 32'b00000000000000000110010111011110; // input=0.650390625, output=0.795847336879
			11'd167: out = 32'b00000000000000000110010110010001; // input=0.654296875, output=0.793476047124
			11'd168: out = 32'b00000000000000000110010101000011; // input=0.658203125, output=0.791092649901
			11'd169: out = 32'b00000000000000000110010011110100; // input=0.662109375, output=0.788697181577
			11'd170: out = 32'b00000000000000000110010010100101; // input=0.666015625, output=0.786289678704
			11'd171: out = 32'b00000000000000000110010001010110; // input=0.669921875, output=0.783870178019
			11'd172: out = 32'b00000000000000000110010000000110; // input=0.673828125, output=0.781438716439
			11'd173: out = 32'b00000000000000000110001110110110; // input=0.677734375, output=0.778995331066
			11'd174: out = 32'b00000000000000000110001101100110; // input=0.681640625, output=0.776540059182
			11'd175: out = 32'b00000000000000000110001100010101; // input=0.685546875, output=0.774072938252
			11'd176: out = 32'b00000000000000000110001011000100; // input=0.689453125, output=0.771594005922
			11'd177: out = 32'b00000000000000000110001001110010; // input=0.693359375, output=0.769103300017
			11'd178: out = 32'b00000000000000000110001000100000; // input=0.697265625, output=0.766600858541
			11'd179: out = 32'b00000000000000000110000111001110; // input=0.701171875, output=0.76408671968
			11'd180: out = 32'b00000000000000000110000101111011; // input=0.705078125, output=0.761560921795
			11'd181: out = 32'b00000000000000000110000100101000; // input=0.708984375, output=0.759023503428
			11'd182: out = 32'b00000000000000000110000011010100; // input=0.712890625, output=0.756474503295
			11'd183: out = 32'b00000000000000000110000010000000; // input=0.716796875, output=0.753913960293
			11'd184: out = 32'b00000000000000000110000000101100; // input=0.720703125, output=0.751341913491
			11'd185: out = 32'b00000000000000000101111111010111; // input=0.724609375, output=0.748758402136
			11'd186: out = 32'b00000000000000000101111110000010; // input=0.728515625, output=0.746163465649
			11'd187: out = 32'b00000000000000000101111100101101; // input=0.732421875, output=0.743557143625
			11'd188: out = 32'b00000000000000000101111011010111; // input=0.736328125, output=0.740939475835
			11'd189: out = 32'b00000000000000000101111010000001; // input=0.740234375, output=0.738310502219
			11'd190: out = 32'b00000000000000000101111000101010; // input=0.744140625, output=0.735670262894
			11'd191: out = 32'b00000000000000000101110111010100; // input=0.748046875, output=0.733018798145
			11'd192: out = 32'b00000000000000000101110101111100; // input=0.751953125, output=0.730356148432
			11'd193: out = 32'b00000000000000000101110100100101; // input=0.755859375, output=0.727682354382
			11'd194: out = 32'b00000000000000000101110011001101; // input=0.759765625, output=0.724997456795
			11'd195: out = 32'b00000000000000000101110001110100; // input=0.763671875, output=0.722301496639
			11'd196: out = 32'b00000000000000000101110000011100; // input=0.767578125, output=0.71959451505
			11'd197: out = 32'b00000000000000000101101111000011; // input=0.771484375, output=0.716876553335
			11'd198: out = 32'b00000000000000000101101101101001; // input=0.775390625, output=0.714147652965
			11'd199: out = 32'b00000000000000000101101100001111; // input=0.779296875, output=0.711407855581
			11'd200: out = 32'b00000000000000000101101010110101; // input=0.783203125, output=0.708657202988
			11'd201: out = 32'b00000000000000000101101001011011; // input=0.787109375, output=0.705895737158
			11'd202: out = 32'b00000000000000000101101000000000; // input=0.791015625, output=0.703123500228
			11'd203: out = 32'b00000000000000000101100110100101; // input=0.794921875, output=0.700340534498
			11'd204: out = 32'b00000000000000000101100101001001; // input=0.798828125, output=0.697546882433
			11'd205: out = 32'b00000000000000000101100011101101; // input=0.802734375, output=0.694742586661
			11'd206: out = 32'b00000000000000000101100010010001; // input=0.806640625, output=0.691927689972
			11'd207: out = 32'b00000000000000000101100000110101; // input=0.810546875, output=0.689102235318
			11'd208: out = 32'b00000000000000000101011111011000; // input=0.814453125, output=0.686266265812
			11'd209: out = 32'b00000000000000000101011101111010; // input=0.818359375, output=0.683419824726
			11'd210: out = 32'b00000000000000000101011100011101; // input=0.822265625, output=0.680562955495
			11'd211: out = 32'b00000000000000000101011010111111; // input=0.826171875, output=0.677695701711
			11'd212: out = 32'b00000000000000000101011001100000; // input=0.830078125, output=0.674818107123
			11'd213: out = 32'b00000000000000000101011000000010; // input=0.833984375, output=0.671930215642
			11'd214: out = 32'b00000000000000000101010110100011; // input=0.837890625, output=0.669032071333
			11'd215: out = 32'b00000000000000000101010101000100; // input=0.841796875, output=0.666123718417
			11'd216: out = 32'b00000000000000000101010011100100; // input=0.845703125, output=0.663205201273
			11'd217: out = 32'b00000000000000000101010010000100; // input=0.849609375, output=0.660276564433
			11'd218: out = 32'b00000000000000000101010000100100; // input=0.853515625, output=0.657337852585
			11'd219: out = 32'b00000000000000000101001111000011; // input=0.857421875, output=0.654389110571
			11'd220: out = 32'b00000000000000000101001101100010; // input=0.861328125, output=0.651430383384
			11'd221: out = 32'b00000000000000000101001100000001; // input=0.865234375, output=0.64846171617
			11'd222: out = 32'b00000000000000000101001010011111; // input=0.869140625, output=0.645483154229
			11'd223: out = 32'b00000000000000000101001000111101; // input=0.873046875, output=0.642494743009
			11'd224: out = 32'b00000000000000000101000111011011; // input=0.876953125, output=0.63949652811
			11'd225: out = 32'b00000000000000000101000101111000; // input=0.880859375, output=0.63648855528
			11'd226: out = 32'b00000000000000000101000100010110; // input=0.884765625, output=0.633470870418
			11'd227: out = 32'b00000000000000000101000010110010; // input=0.888671875, output=0.63044351957
			11'd228: out = 32'b00000000000000000101000001001111; // input=0.892578125, output=0.62740654893
			11'd229: out = 32'b00000000000000000100111111101011; // input=0.896484375, output=0.624360004837
			11'd230: out = 32'b00000000000000000100111110000111; // input=0.900390625, output=0.621303933779
			11'd231: out = 32'b00000000000000000100111100100010; // input=0.904296875, output=0.618238382388
			11'd232: out = 32'b00000000000000000100111010111110; // input=0.908203125, output=0.615163397439
			11'd233: out = 32'b00000000000000000100111001011001; // input=0.912109375, output=0.612079025854
			11'd234: out = 32'b00000000000000000100110111110011; // input=0.916015625, output=0.608985314696
			11'd235: out = 32'b00000000000000000100110110001110; // input=0.919921875, output=0.605882311171
			11'd236: out = 32'b00000000000000000100110100101000; // input=0.923828125, output=0.602770062628
			11'd237: out = 32'b00000000000000000100110011000001; // input=0.927734375, output=0.599648616555
			11'd238: out = 32'b00000000000000000100110001011011; // input=0.931640625, output=0.596518020582
			11'd239: out = 32'b00000000000000000100101111110100; // input=0.935546875, output=0.593378322478
			11'd240: out = 32'b00000000000000000100101110001101; // input=0.939453125, output=0.590229570151
			11'd241: out = 32'b00000000000000000100101100100101; // input=0.943359375, output=0.587071811646
			11'd242: out = 32'b00000000000000000100101010111101; // input=0.947265625, output=0.583905095149
			11'd243: out = 32'b00000000000000000100101001010101; // input=0.951171875, output=0.580729468977
			11'd244: out = 32'b00000000000000000100100111101101; // input=0.955078125, output=0.577544981589
			11'd245: out = 32'b00000000000000000100100110000100; // input=0.958984375, output=0.574351681575
			11'd246: out = 32'b00000000000000000100100100011011; // input=0.962890625, output=0.571149617661
			11'd247: out = 32'b00000000000000000100100010110010; // input=0.966796875, output=0.567938838706
			11'd248: out = 32'b00000000000000000100100001001001; // input=0.970703125, output=0.564719393703
			11'd249: out = 32'b00000000000000000100011111011111; // input=0.974609375, output=0.561491331777
			11'd250: out = 32'b00000000000000000100011101110101; // input=0.978515625, output=0.558254702185
			11'd251: out = 32'b00000000000000000100011100001011; // input=0.982421875, output=0.555009554312
			11'd252: out = 32'b00000000000000000100011010100000; // input=0.986328125, output=0.551755937677
			11'd253: out = 32'b00000000000000000100011000110101; // input=0.990234375, output=0.548493901924
			11'd254: out = 32'b00000000000000000100010111001010; // input=0.994140625, output=0.54522349683
			11'd255: out = 32'b00000000000000000100010101011110; // input=0.998046875, output=0.541944772296
			11'd256: out = 32'b00000000000000000100010011110011; // input=1.001953125, output=0.538657778351
			11'd257: out = 32'b00000000000000000100010010000111; // input=1.005859375, output=0.535362565152
			11'd258: out = 32'b00000000000000000100010000011011; // input=1.009765625, output=0.532059182978
			11'd259: out = 32'b00000000000000000100001110101110; // input=1.013671875, output=0.528747682236
			11'd260: out = 32'b00000000000000000100001101000001; // input=1.017578125, output=0.525428113455
			11'd261: out = 32'b00000000000000000100001011010100; // input=1.021484375, output=0.522100527287
			11'd262: out = 32'b00000000000000000100001001100111; // input=1.025390625, output=0.518764974507
			11'd263: out = 32'b00000000000000000100000111111001; // input=1.029296875, output=0.515421506013
			11'd264: out = 32'b00000000000000000100000110001100; // input=1.033203125, output=0.51207017282
			11'd265: out = 32'b00000000000000000100000100011101; // input=1.037109375, output=0.508711026066
			11'd266: out = 32'b00000000000000000100000010101111; // input=1.041015625, output=0.505344117008
			11'd267: out = 32'b00000000000000000100000001000001; // input=1.044921875, output=0.501969497021
			11'd268: out = 32'b00000000000000000011111111010010; // input=1.048828125, output=0.498587217597
			11'd269: out = 32'b00000000000000000011111101100011; // input=1.052734375, output=0.495197330345
			11'd270: out = 32'b00000000000000000011111011110011; // input=1.056640625, output=0.491799886991
			11'd271: out = 32'b00000000000000000011111010000100; // input=1.060546875, output=0.488394939376
			11'd272: out = 32'b00000000000000000011111000010100; // input=1.064453125, output=0.484982539455
			11'd273: out = 32'b00000000000000000011110110100100; // input=1.068359375, output=0.481562739297
			11'd274: out = 32'b00000000000000000011110100110100; // input=1.072265625, output=0.478135591084
			11'd275: out = 32'b00000000000000000011110011000011; // input=1.076171875, output=0.474701147111
			11'd276: out = 32'b00000000000000000011110001010010; // input=1.080078125, output=0.471259459782
			11'd277: out = 32'b00000000000000000011101111100001; // input=1.083984375, output=0.467810581613
			11'd278: out = 32'b00000000000000000011101101110000; // input=1.087890625, output=0.464354565231
			11'd279: out = 32'b00000000000000000011101011111110; // input=1.091796875, output=0.460891463369
			11'd280: out = 32'b00000000000000000011101010001101; // input=1.095703125, output=0.45742132887
			11'd281: out = 32'b00000000000000000011101000011011; // input=1.099609375, output=0.453944214685
			11'd282: out = 32'b00000000000000000011100110101001; // input=1.103515625, output=0.45046017387
			11'd283: out = 32'b00000000000000000011100100110110; // input=1.107421875, output=0.446969259586
			11'd284: out = 32'b00000000000000000011100011000100; // input=1.111328125, output=0.443471525102
			11'd285: out = 32'b00000000000000000011100001010001; // input=1.115234375, output=0.439967023787
			11'd286: out = 32'b00000000000000000011011111011110; // input=1.119140625, output=0.436455809118
			11'd287: out = 32'b00000000000000000011011101101011; // input=1.123046875, output=0.432937934669
			11'd288: out = 32'b00000000000000000011011011110111; // input=1.126953125, output=0.429413454121
			11'd289: out = 32'b00000000000000000011011010000011; // input=1.130859375, output=0.425882421251
			11'd290: out = 32'b00000000000000000011011000001111; // input=1.134765625, output=0.42234488994
			11'd291: out = 32'b00000000000000000011010110011011; // input=1.138671875, output=0.418800914165
			11'd292: out = 32'b00000000000000000011010100100111; // input=1.142578125, output=0.415250548003
			11'd293: out = 32'b00000000000000000011010010110010; // input=1.146484375, output=0.411693845629
			11'd294: out = 32'b00000000000000000011010000111110; // input=1.150390625, output=0.408130861314
			11'd295: out = 32'b00000000000000000011001111001001; // input=1.154296875, output=0.404561649424
			11'd296: out = 32'b00000000000000000011001101010100; // input=1.158203125, output=0.40098626442
			11'd297: out = 32'b00000000000000000011001011011110; // input=1.162109375, output=0.39740476086
			11'd298: out = 32'b00000000000000000011001001101001; // input=1.166015625, output=0.393817193392
			11'd299: out = 32'b00000000000000000011000111110011; // input=1.169921875, output=0.390223616758
			11'd300: out = 32'b00000000000000000011000101111101; // input=1.173828125, output=0.386624085792
			11'd301: out = 32'b00000000000000000011000100000111; // input=1.177734375, output=0.383018655418
			11'd302: out = 32'b00000000000000000011000010010000; // input=1.181640625, output=0.37940738065
			11'd303: out = 32'b00000000000000000011000000011010; // input=1.185546875, output=0.375790316593
			11'd304: out = 32'b00000000000000000010111110100011; // input=1.189453125, output=0.372167518438
			11'd305: out = 32'b00000000000000000010111100101100; // input=1.193359375, output=0.368539041464
			11'd306: out = 32'b00000000000000000010111010110101; // input=1.197265625, output=0.364904941038
			11'd307: out = 32'b00000000000000000010111000111110; // input=1.201171875, output=0.361265272612
			11'd308: out = 32'b00000000000000000010110111000110; // input=1.205078125, output=0.357620091721
			11'd309: out = 32'b00000000000000000010110101001111; // input=1.208984375, output=0.353969453989
			11'd310: out = 32'b00000000000000000010110011010111; // input=1.212890625, output=0.350313415118
			11'd311: out = 32'b00000000000000000010110001011111; // input=1.216796875, output=0.346652030895
			11'd312: out = 32'b00000000000000000010101111100111; // input=1.220703125, output=0.342985357189
			11'd313: out = 32'b00000000000000000010101101101111; // input=1.224609375, output=0.339313449948
			11'd314: out = 32'b00000000000000000010101011110110; // input=1.228515625, output=0.335636365202
			11'd315: out = 32'b00000000000000000010101001111101; // input=1.232421875, output=0.331954159057
			11'd316: out = 32'b00000000000000000010101000000101; // input=1.236328125, output=0.328266887701
			11'd317: out = 32'b00000000000000000010100110001100; // input=1.240234375, output=0.324574607395
			11'd318: out = 32'b00000000000000000010100100010011; // input=1.244140625, output=0.320877374481
			11'd319: out = 32'b00000000000000000010100010011001; // input=1.248046875, output=0.317175245372
			11'd320: out = 32'b00000000000000000010100000100000; // input=1.251953125, output=0.31346827656
			11'd321: out = 32'b00000000000000000010011110100110; // input=1.255859375, output=0.309756524607
			11'd322: out = 32'b00000000000000000010011100101100; // input=1.259765625, output=0.306040046151
			11'd323: out = 32'b00000000000000000010011010110010; // input=1.263671875, output=0.3023188979
			11'd324: out = 32'b00000000000000000010011000111000; // input=1.267578125, output=0.298593136635
			11'd325: out = 32'b00000000000000000010010110111110; // input=1.271484375, output=0.294862819205
			11'd326: out = 32'b00000000000000000010010101000100; // input=1.275390625, output=0.291128002532
			11'd327: out = 32'b00000000000000000010010011001001; // input=1.279296875, output=0.287388743604
			11'd328: out = 32'b00000000000000000010010001001110; // input=1.283203125, output=0.283645099478
			11'd329: out = 32'b00000000000000000010001111010100; // input=1.287109375, output=0.279897127276
			11'd330: out = 32'b00000000000000000010001101011001; // input=1.291015625, output=0.276144884188
			11'd331: out = 32'b00000000000000000010001011011110; // input=1.294921875, output=0.272388427469
			11'd332: out = 32'b00000000000000000010001001100010; // input=1.298828125, output=0.268627814438
			11'd333: out = 32'b00000000000000000010000111100111; // input=1.302734375, output=0.264863102477
			11'd334: out = 32'b00000000000000000010000101101100; // input=1.306640625, output=0.26109434903
			11'd335: out = 32'b00000000000000000010000011110000; // input=1.310546875, output=0.257321611606
			11'd336: out = 32'b00000000000000000010000001110100; // input=1.314453125, output=0.25354494777
			11'd337: out = 32'b00000000000000000001111111111000; // input=1.318359375, output=0.24976441515
			11'd338: out = 32'b00000000000000000001111101111100; // input=1.322265625, output=0.245980071432
			11'd339: out = 32'b00000000000000000001111100000000; // input=1.326171875, output=0.242191974361
			11'd340: out = 32'b00000000000000000001111010000100; // input=1.330078125, output=0.238400181739
			11'd341: out = 32'b00000000000000000001111000001000; // input=1.333984375, output=0.234604751423
			11'd342: out = 32'b00000000000000000001110110001011; // input=1.337890625, output=0.230805741327
			11'd343: out = 32'b00000000000000000001110100001110; // input=1.341796875, output=0.22700320942
			11'd344: out = 32'b00000000000000000001110010010010; // input=1.345703125, output=0.223197213723
			11'd345: out = 32'b00000000000000000001110000010101; // input=1.349609375, output=0.219387812311
			11'd346: out = 32'b00000000000000000001101110011000; // input=1.353515625, output=0.215575063311
			11'd347: out = 32'b00000000000000000001101100011011; // input=1.357421875, output=0.211759024901
			11'd348: out = 32'b00000000000000000001101010011110; // input=1.361328125, output=0.207939755308
			11'd349: out = 32'b00000000000000000001101000100001; // input=1.365234375, output=0.204117312811
			11'd350: out = 32'b00000000000000000001100110100011; // input=1.369140625, output=0.200291755735
			11'd351: out = 32'b00000000000000000001100100100110; // input=1.373046875, output=0.196463142453
			11'd352: out = 32'b00000000000000000001100010101000; // input=1.376953125, output=0.192631531385
			11'd353: out = 32'b00000000000000000001100000101010; // input=1.380859375, output=0.188796980997
			11'd354: out = 32'b00000000000000000001011110101101; // input=1.384765625, output=0.184959549799
			11'd355: out = 32'b00000000000000000001011100101111; // input=1.388671875, output=0.181119296346
			11'd356: out = 32'b00000000000000000001011010110001; // input=1.392578125, output=0.177276279236
			11'd357: out = 32'b00000000000000000001011000110011; // input=1.396484375, output=0.173430557107
			11'd358: out = 32'b00000000000000000001010110110101; // input=1.400390625, output=0.169582188642
			11'd359: out = 32'b00000000000000000001010100110111; // input=1.404296875, output=0.165731232561
			11'd360: out = 32'b00000000000000000001010010111000; // input=1.408203125, output=0.161877747625
			11'd361: out = 32'b00000000000000000001010000111010; // input=1.412109375, output=0.158021792634
			11'd362: out = 32'b00000000000000000001001110111100; // input=1.416015625, output=0.154163426425
			11'd363: out = 32'b00000000000000000001001100111101; // input=1.419921875, output=0.150302707872
			11'd364: out = 32'b00000000000000000001001010111111; // input=1.423828125, output=0.146439695884
			11'd365: out = 32'b00000000000000000001001001000000; // input=1.427734375, output=0.142574449407
			11'd366: out = 32'b00000000000000000001000111000001; // input=1.431640625, output=0.138707027419
			11'd367: out = 32'b00000000000000000001000101000010; // input=1.435546875, output=0.134837488933
			11'd368: out = 32'b00000000000000000001000011000011; // input=1.439453125, output=0.130965892992
			11'd369: out = 32'b00000000000000000001000001000101; // input=1.443359375, output=0.127092298673
			11'd370: out = 32'b00000000000000000000111111000110; // input=1.447265625, output=0.123216765082
			11'd371: out = 32'b00000000000000000000111101000111; // input=1.451171875, output=0.119339351355
			11'd372: out = 32'b00000000000000000000111011000111; // input=1.455078125, output=0.115460116656
			11'd373: out = 32'b00000000000000000000111001001000; // input=1.458984375, output=0.111579120177
			11'd374: out = 32'b00000000000000000000110111001001; // input=1.462890625, output=0.107696421139
			11'd375: out = 32'b00000000000000000000110101001010; // input=1.466796875, output=0.103812078785
			11'd376: out = 32'b00000000000000000000110011001010; // input=1.470703125, output=0.0999261523872
			11'd377: out = 32'b00000000000000000000110001001011; // input=1.474609375, output=0.0960387012391
			11'd378: out = 32'b00000000000000000000101111001100; // input=1.478515625, output=0.0921497846586
			11'd379: out = 32'b00000000000000000000101101001100; // input=1.482421875, output=0.0882594619857
			11'd380: out = 32'b00000000000000000000101011001101; // input=1.486328125, output=0.084367792582
			11'd381: out = 32'b00000000000000000000101001001101; // input=1.490234375, output=0.0804748358296
			11'd382: out = 32'b00000000000000000000100111001101; // input=1.494140625, output=0.0765806511302
			11'd383: out = 32'b00000000000000000000100101001110; // input=1.498046875, output=0.0726852979043
			11'd384: out = 32'b00000000000000000000100011001110; // input=1.501953125, output=0.0687888355902
			11'd385: out = 32'b00000000000000000000100001001110; // input=1.505859375, output=0.0648913236431
			11'd386: out = 32'b00000000000000000000011111001111; // input=1.509765625, output=0.0609928215342
			11'd387: out = 32'b00000000000000000000011101001111; // input=1.513671875, output=0.0570933887499
			11'd388: out = 32'b00000000000000000000011011001111; // input=1.517578125, output=0.0531930847907
			11'd389: out = 32'b00000000000000000000011001001111; // input=1.521484375, output=0.0492919691706
			11'd390: out = 32'b00000000000000000000010111001111; // input=1.525390625, output=0.0453901014156
			11'd391: out = 32'b00000000000000000000010101001111; // input=1.529296875, output=0.0414875410635
			11'd392: out = 32'b00000000000000000000010011010000; // input=1.533203125, output=0.0375843476626
			11'd393: out = 32'b00000000000000000000010001010000; // input=1.537109375, output=0.0336805807707
			11'd394: out = 32'b00000000000000000000001111010000; // input=1.541015625, output=0.0297762999547
			11'd395: out = 32'b00000000000000000000001101010000; // input=1.544921875, output=0.0258715647889
			11'd396: out = 32'b00000000000000000000001011010000; // input=1.548828125, output=0.0219664348549
			11'd397: out = 32'b00000000000000000000001001010000; // input=1.552734375, output=0.0180609697401
			11'd398: out = 32'b00000000000000000000000111010000; // input=1.556640625, output=0.0141552290372
			11'd399: out = 32'b00000000000000000000000101010000; // input=1.560546875, output=0.0102492723429
			11'd400: out = 32'b00000000000000000000000011010000; // input=1.564453125, output=0.00634315925725
			11'd401: out = 32'b00000000000000000000000001010000; // input=1.568359375, output=0.00243694938283
			11'd402: out = 32'b10000000000000000000000000110000; // input=1.572265625, output=-0.00146929767644
			11'd403: out = 32'b10000000000000000000000010110000; // input=1.576171875, output=-0.00537552231604
			11'd404: out = 32'b10000000000000000000000100110000; // input=1.580078125, output=-0.00928166493177
			11'd405: out = 32'b10000000000000000000000110110000; // input=1.583984375, output=-0.0131876659207
			11'd406: out = 32'b10000000000000000000001000110000; // input=1.587890625, output=-0.0170934656821
			11'd407: out = 32'b10000000000000000000001010110000; // input=1.591796875, output=-0.0209990046183
			11'd408: out = 32'b10000000000000000000001100110000; // input=1.595703125, output=-0.0249042231354
			11'd409: out = 32'b10000000000000000000001110110000; // input=1.599609375, output=-0.0288090616448
			11'd410: out = 32'b10000000000000000000010000110000; // input=1.603515625, output=-0.0327134605633
			11'd411: out = 32'b10000000000000000000010010110000; // input=1.607421875, output=-0.0366173603147
			11'd412: out = 32'b10000000000000000000010100110000; // input=1.611328125, output=-0.0405207013302
			11'd413: out = 32'b10000000000000000000010110110000; // input=1.615234375, output=-0.0444234240496
			11'd414: out = 32'b10000000000000000000011000110000; // input=1.619140625, output=-0.0483254689223
			11'd415: out = 32'b10000000000000000000011010101111; // input=1.623046875, output=-0.0522267764077
			11'd416: out = 32'b10000000000000000000011100101111; // input=1.626953125, output=-0.0561272869768
			11'd417: out = 32'b10000000000000000000011110101111; // input=1.630859375, output=-0.0600269411126
			11'd418: out = 32'b10000000000000000000100000101111; // input=1.634765625, output=-0.0639256793111
			11'd419: out = 32'b10000000000000000000100010101110; // input=1.638671875, output=-0.0678234420824
			11'd420: out = 32'b10000000000000000000100100101110; // input=1.642578125, output=-0.0717201699514
			11'd421: out = 32'b10000000000000000000100110101110; // input=1.646484375, output=-0.0756158034588
			11'd422: out = 32'b10000000000000000000101000101101; // input=1.650390625, output=-0.0795102831621
			11'd423: out = 32'b10000000000000000000101010101101; // input=1.654296875, output=-0.0834035496363
			11'd424: out = 32'b10000000000000000000101100101101; // input=1.658203125, output=-0.087295543475
			11'd425: out = 32'b10000000000000000000101110101100; // input=1.662109375, output=-0.0911862052911
			11'd426: out = 32'b10000000000000000000110000101011; // input=1.666015625, output=-0.0950754757179
			11'd427: out = 32'b10000000000000000000110010101011; // input=1.669921875, output=-0.0989632954099
			11'd428: out = 32'b10000000000000000000110100101010; // input=1.673828125, output=-0.102849605044
			11'd429: out = 32'b10000000000000000000110110101001; // input=1.677734375, output=-0.106734345319
			11'd430: out = 32'b10000000000000000000111000101001; // input=1.681640625, output=-0.11061745696
			11'd431: out = 32'b10000000000000000000111010101000; // input=1.685546875, output=-0.114498880714
			11'd432: out = 32'b10000000000000000000111100100111; // input=1.689453125, output=-0.118378557356
			11'd433: out = 32'b10000000000000000000111110100110; // input=1.693359375, output=-0.122256427688
			11'd434: out = 32'b10000000000000000001000000100101; // input=1.697265625, output=-0.126132432536
			11'd435: out = 32'b10000000000000000001000010100100; // input=1.701171875, output=-0.130006512759
			11'd436: out = 32'b10000000000000000001000100100011; // input=1.705078125, output=-0.133878609242
			11'd437: out = 32'b10000000000000000001000110100010; // input=1.708984375, output=-0.137748662903
			11'd438: out = 32'b10000000000000000001001000100000; // input=1.712890625, output=-0.141616614688
			11'd439: out = 32'b10000000000000000001001010011111; // input=1.716796875, output=-0.145482405578
			11'd440: out = 32'b10000000000000000001001100011110; // input=1.720703125, output=-0.149345976585
			11'd441: out = 32'b10000000000000000001001110011100; // input=1.724609375, output=-0.153207268757
			11'd442: out = 32'b10000000000000000001010000011011; // input=1.728515625, output=-0.157066223174
			11'd443: out = 32'b10000000000000000001010010011001; // input=1.732421875, output=-0.160922780954
			11'd444: out = 32'b10000000000000000001010100010111; // input=1.736328125, output=-0.164776883251
			11'd445: out = 32'b10000000000000000001010110010110; // input=1.740234375, output=-0.168628471254
			11'd446: out = 32'b10000000000000000001011000010100; // input=1.744140625, output=-0.172477486195
			11'd447: out = 32'b10000000000000000001011010010010; // input=1.748046875, output=-0.176323869342
			11'd448: out = 32'b10000000000000000001011100010000; // input=1.751953125, output=-0.180167562003
			11'd449: out = 32'b10000000000000000001011110001110; // input=1.755859375, output=-0.184008505529
			11'd450: out = 32'b10000000000000000001100000001011; // input=1.759765625, output=-0.187846641311
			11'd451: out = 32'b10000000000000000001100010001001; // input=1.763671875, output=-0.191681910785
			11'd452: out = 32'b10000000000000000001100100000111; // input=1.767578125, output=-0.195514255429
			11'd453: out = 32'b10000000000000000001100110000100; // input=1.771484375, output=-0.199343616766
			11'd454: out = 32'b10000000000000000001101000000001; // input=1.775390625, output=-0.203169936364
			11'd455: out = 32'b10000000000000000001101001111111; // input=1.779296875, output=-0.206993155839
			11'd456: out = 32'b10000000000000000001101011111100; // input=1.783203125, output=-0.210813216853
			11'd457: out = 32'b10000000000000000001101101111001; // input=1.787109375, output=-0.214630061117
			11'd458: out = 32'b10000000000000000001101111110110; // input=1.791015625, output=-0.218443630391
			11'd459: out = 32'b10000000000000000001110001110011; // input=1.794921875, output=-0.222253866483
			11'd460: out = 32'b10000000000000000001110011110000; // input=1.798828125, output=-0.226060711255
			11'd461: out = 32'b10000000000000000001110101101100; // input=1.802734375, output=-0.229864106618
			11'd462: out = 32'b10000000000000000001110111101001; // input=1.806640625, output=-0.233663994538
			11'd463: out = 32'b10000000000000000001111001100101; // input=1.810546875, output=-0.237460317033
			11'd464: out = 32'b10000000000000000001111011100001; // input=1.814453125, output=-0.241253016175
			11'd465: out = 32'b10000000000000000001111101011110; // input=1.818359375, output=-0.245042034094
			11'd466: out = 32'b10000000000000000001111111011010; // input=1.822265625, output=-0.248827312972
			11'd467: out = 32'b10000000000000000010000001010101; // input=1.826171875, output=-0.252608795052
			11'd468: out = 32'b10000000000000000010000011010001; // input=1.830078125, output=-0.256386422632
			11'd469: out = 32'b10000000000000000010000101001101; // input=1.833984375, output=-0.260160138071
			11'd470: out = 32'b10000000000000000010000111001000; // input=1.837890625, output=-0.263929883786
			11'd471: out = 32'b10000000000000000010001001000100; // input=1.841796875, output=-0.267695602256
			11'd472: out = 32'b10000000000000000010001010111111; // input=1.845703125, output=-0.271457236021
			11'd473: out = 32'b10000000000000000010001100111010; // input=1.849609375, output=-0.275214727682
			11'd474: out = 32'b10000000000000000010001110110101; // input=1.853515625, output=-0.278968019905
			11'd475: out = 32'b10000000000000000010010000110000; // input=1.857421875, output=-0.282717055419
			11'd476: out = 32'b10000000000000000010010010101011; // input=1.861328125, output=-0.286461777019
			11'd477: out = 32'b10000000000000000010010100100101; // input=1.865234375, output=-0.290202127564
			11'd478: out = 32'b10000000000000000010010110100000; // input=1.869140625, output=-0.293938049982
			11'd479: out = 32'b10000000000000000010011000011010; // input=1.873046875, output=-0.297669487267
			11'd480: out = 32'b10000000000000000010011010010100; // input=1.876953125, output=-0.301396382482
			11'd481: out = 32'b10000000000000000010011100001110; // input=1.880859375, output=-0.305118678759
			11'd482: out = 32'b10000000000000000010011110001000; // input=1.884765625, output=-0.308836319301
			11'd483: out = 32'b10000000000000000010100000000010; // input=1.888671875, output=-0.31254924738
			11'd484: out = 32'b10000000000000000010100001111011; // input=1.892578125, output=-0.316257406342
			11'd485: out = 32'b10000000000000000010100011110100; // input=1.896484375, output=-0.319960739605
			11'd486: out = 32'b10000000000000000010100101101110; // input=1.900390625, output=-0.323659190661
			11'd487: out = 32'b10000000000000000010100111100111; // input=1.904296875, output=-0.327352703076
			11'd488: out = 32'b10000000000000000010101001100000; // input=1.908203125, output=-0.331041220491
			11'd489: out = 32'b10000000000000000010101011011000; // input=1.912109375, output=-0.334724686625
			11'd490: out = 32'b10000000000000000010101101010001; // input=1.916015625, output=-0.338403045272
			11'd491: out = 32'b10000000000000000010101111001001; // input=1.919921875, output=-0.342076240304
			11'd492: out = 32'b10000000000000000010110001000001; // input=1.923828125, output=-0.345744215674
			11'd493: out = 32'b10000000000000000010110010111001; // input=1.927734375, output=-0.349406915413
			11'd494: out = 32'b10000000000000000010110100110001; // input=1.931640625, output=-0.353064283632
			11'd495: out = 32'b10000000000000000010110110101001; // input=1.935546875, output=-0.356716264525
			11'd496: out = 32'b10000000000000000010111000100000; // input=1.939453125, output=-0.360362802366
			11'd497: out = 32'b10000000000000000010111010011000; // input=1.943359375, output=-0.364003841514
			11'd498: out = 32'b10000000000000000010111100001111; // input=1.947265625, output=-0.367639326412
			11'd499: out = 32'b10000000000000000010111110000110; // input=1.951171875, output=-0.371269201585
			11'd500: out = 32'b10000000000000000010111111111101; // input=1.955078125, output=-0.374893411648
			11'd501: out = 32'b10000000000000000011000001110011; // input=1.958984375, output=-0.378511901298
			11'd502: out = 32'b10000000000000000011000011101001; // input=1.962890625, output=-0.382124615322
			11'd503: out = 32'b10000000000000000011000101100000; // input=1.966796875, output=-0.385731498595
			11'd504: out = 32'b10000000000000000011000111010110; // input=1.970703125, output=-0.38933249608
			11'd505: out = 32'b10000000000000000011001001001011; // input=1.974609375, output=-0.392927552829
			11'd506: out = 32'b10000000000000000011001011000001; // input=1.978515625, output=-0.396516613988
			11'd507: out = 32'b10000000000000000011001100110110; // input=1.982421875, output=-0.400099624791
			11'd508: out = 32'b10000000000000000011001110101100; // input=1.986328125, output=-0.403676530566
			11'd509: out = 32'b10000000000000000011010000100001; // input=1.990234375, output=-0.407247276734
			11'd510: out = 32'b10000000000000000011010010010101; // input=1.994140625, output=-0.41081180881
			11'd511: out = 32'b10000000000000000011010100001010; // input=1.998046875, output=-0.414370072403
			11'd512: out = 32'b10000000000000000011010101111110; // input=2.001953125, output=-0.417922013218
			11'd513: out = 32'b10000000000000000011010111110011; // input=2.005859375, output=-0.421467577057
			11'd514: out = 32'b10000000000000000011011001100111; // input=2.009765625, output=-0.42500670982
			11'd515: out = 32'b10000000000000000011011011011010; // input=2.013671875, output=-0.428539357504
			11'd516: out = 32'b10000000000000000011011101001110; // input=2.017578125, output=-0.432065466204
			11'd517: out = 32'b10000000000000000011011111000001; // input=2.021484375, output=-0.435584982116
			11'd518: out = 32'b10000000000000000011100000110100; // input=2.025390625, output=-0.439097851538
			11'd519: out = 32'b10000000000000000011100010100111; // input=2.029296875, output=-0.442604020867
			11'd520: out = 32'b10000000000000000011100100011010; // input=2.033203125, output=-0.446103436603
			11'd521: out = 32'b10000000000000000011100110001100; // input=2.037109375, output=-0.449596045349
			11'd522: out = 32'b10000000000000000011100111111111; // input=2.041015625, output=-0.453081793813
			11'd523: out = 32'b10000000000000000011101001110001; // input=2.044921875, output=-0.456560628806
			11'd524: out = 32'b10000000000000000011101011100010; // input=2.048828125, output=-0.460032497246
			11'd525: out = 32'b10000000000000000011101101010100; // input=2.052734375, output=-0.463497346155
			11'd526: out = 32'b10000000000000000011101111000101; // input=2.056640625, output=-0.466955122666
			11'd527: out = 32'b10000000000000000011110000110110; // input=2.060546875, output=-0.470405774016
			11'd528: out = 32'b10000000000000000011110010100111; // input=2.064453125, output=-0.473849247552
			11'd529: out = 32'b10000000000000000011110100011000; // input=2.068359375, output=-0.477285490732
			11'd530: out = 32'b10000000000000000011110110001000; // input=2.072265625, output=-0.480714451123
			11'd531: out = 32'b10000000000000000011110111111000; // input=2.076171875, output=-0.484136076402
			11'd532: out = 32'b10000000000000000011111001101000; // input=2.080078125, output=-0.487550314361
			11'd533: out = 32'b10000000000000000011111011011000; // input=2.083984375, output=-0.490957112901
			11'd534: out = 32'b10000000000000000011111101000111; // input=2.087890625, output=-0.49435642004
			11'd535: out = 32'b10000000000000000011111110110110; // input=2.091796875, output=-0.497748183909
			11'd536: out = 32'b10000000000000000100000000100101; // input=2.095703125, output=-0.501132352752
			11'd537: out = 32'b10000000000000000100000010010100; // input=2.099609375, output=-0.504508874933
			11'd538: out = 32'b10000000000000000100000100000010; // input=2.103515625, output=-0.507877698929
			11'd539: out = 32'b10000000000000000100000101110000; // input=2.107421875, output=-0.511238773335
			11'd540: out = 32'b10000000000000000100000111011110; // input=2.111328125, output=-0.514592046868
			11'd541: out = 32'b10000000000000000100001001001100; // input=2.115234375, output=-0.517937468358
			11'd542: out = 32'b10000000000000000100001010111001; // input=2.119140625, output=-0.52127498676
			11'd543: out = 32'b10000000000000000100001100100110; // input=2.123046875, output=-0.524604551148
			11'd544: out = 32'b10000000000000000100001110010011; // input=2.126953125, output=-0.527926110715
			11'd545: out = 32'b10000000000000000100010000000000; // input=2.130859375, output=-0.531239614779
			11'd546: out = 32'b10000000000000000100010001101100; // input=2.134765625, output=-0.53454501278
			11'd547: out = 32'b10000000000000000100010011011000; // input=2.138671875, output=-0.537842254283
			11'd548: out = 32'b10000000000000000100010101000100; // input=2.142578125, output=-0.541131288974
			11'd549: out = 32'b10000000000000000100010110101111; // input=2.146484375, output=-0.544412066667
			11'd550: out = 32'b10000000000000000100011000011011; // input=2.150390625, output=-0.547684537302
			11'd551: out = 32'b10000000000000000100011010000101; // input=2.154296875, output=-0.550948650945
			11'd552: out = 32'b10000000000000000100011011110000; // input=2.158203125, output=-0.554204357789
			11'd553: out = 32'b10000000000000000100011101011011; // input=2.162109375, output=-0.557451608157
			11'd554: out = 32'b10000000000000000100011111000101; // input=2.166015625, output=-0.560690352499
			11'd555: out = 32'b10000000000000000100100000101111; // input=2.169921875, output=-0.563920541396
			11'd556: out = 32'b10000000000000000100100010011000; // input=2.173828125, output=-0.567142125559
			11'd557: out = 32'b10000000000000000100100100000001; // input=2.177734375, output=-0.570355055831
			11'd558: out = 32'b10000000000000000100100101101010; // input=2.181640625, output=-0.573559283187
			11'd559: out = 32'b10000000000000000100100111010011; // input=2.185546875, output=-0.576754758734
			11'd560: out = 32'b10000000000000000100101000111100; // input=2.189453125, output=-0.579941433713
			11'd561: out = 32'b10000000000000000100101010100100; // input=2.193359375, output=-0.583119259499
			11'd562: out = 32'b10000000000000000100101100001011; // input=2.197265625, output=-0.586288187603
			11'd563: out = 32'b10000000000000000100101101110011; // input=2.201171875, output=-0.58944816967
			11'd564: out = 32'b10000000000000000100101111011010; // input=2.205078125, output=-0.592599157484
			11'd565: out = 32'b10000000000000000100110001000001; // input=2.208984375, output=-0.595741102963
			11'd566: out = 32'b10000000000000000100110010101000; // input=2.212890625, output=-0.598873958166
			11'd567: out = 32'b10000000000000000100110100001110; // input=2.216796875, output=-0.601997675289
			11'd568: out = 32'b10000000000000000100110101110100; // input=2.220703125, output=-0.605112206669
			11'd569: out = 32'b10000000000000000100110111011010; // input=2.224609375, output=-0.60821750478
			11'd570: out = 32'b10000000000000000100111001000000; // input=2.228515625, output=-0.611313522241
			11'd571: out = 32'b10000000000000000100111010100101; // input=2.232421875, output=-0.61440021181
			11'd572: out = 32'b10000000000000000100111100001010; // input=2.236328125, output=-0.617477526387
			11'd573: out = 32'b10000000000000000100111101101110; // input=2.240234375, output=-0.620545419017
			11'd574: out = 32'b10000000000000000100111111010010; // input=2.244140625, output=-0.623603842888
			11'd575: out = 32'b10000000000000000101000000110110; // input=2.248046875, output=-0.626652751331
			11'd576: out = 32'b10000000000000000101000010011010; // input=2.251953125, output=-0.629692097824
			11'd577: out = 32'b10000000000000000101000011111101; // input=2.255859375, output=-0.63272183599
			11'd578: out = 32'b10000000000000000101000101100000; // input=2.259765625, output=-0.635741919599
			11'd579: out = 32'b10000000000000000101000111000011; // input=2.263671875, output=-0.638752302569
			11'd580: out = 32'b10000000000000000101001000100101; // input=2.267578125, output=-0.641752938965
			11'd581: out = 32'b10000000000000000101001010000111; // input=2.271484375, output=-0.644743783001
			11'd582: out = 32'b10000000000000000101001011101001; // input=2.275390625, output=-0.647724789039
			11'd583: out = 32'b10000000000000000101001101001010; // input=2.279296875, output=-0.650695911595
			11'd584: out = 32'b10000000000000000101001110101011; // input=2.283203125, output=-0.653657105331
			11'd585: out = 32'b10000000000000000101010000001100; // input=2.287109375, output=-0.656608325064
			11'd586: out = 32'b10000000000000000101010001101100; // input=2.291015625, output=-0.659549525762
			11'd587: out = 32'b10000000000000000101010011001100; // input=2.294921875, output=-0.662480662545
			11'd588: out = 32'b10000000000000000101010100101100; // input=2.298828125, output=-0.665401690689
			11'd589: out = 32'b10000000000000000101010110001011; // input=2.302734375, output=-0.668312565622
			11'd590: out = 32'b10000000000000000101010111101010; // input=2.306640625, output=-0.671213242927
			11'd591: out = 32'b10000000000000000101011001001001; // input=2.310546875, output=-0.674103678343
			11'd592: out = 32'b10000000000000000101011010100111; // input=2.314453125, output=-0.676983827767
			11'd593: out = 32'b10000000000000000101011100000101; // input=2.318359375, output=-0.679853647251
			11'd594: out = 32'b10000000000000000101011101100011; // input=2.322265625, output=-0.682713093005
			11'd595: out = 32'b10000000000000000101011111000000; // input=2.326171875, output=-0.685562121397
			11'd596: out = 32'b10000000000000000101100000011110; // input=2.330078125, output=-0.688400688954
			11'd597: out = 32'b10000000000000000101100001111010; // input=2.333984375, output=-0.691228752363
			11'd598: out = 32'b10000000000000000101100011010111; // input=2.337890625, output=-0.694046268473
			11'd599: out = 32'b10000000000000000101100100110010; // input=2.341796875, output=-0.69685319429
			11'd600: out = 32'b10000000000000000101100110001110; // input=2.345703125, output=-0.699649486985
			11'd601: out = 32'b10000000000000000101100111101001; // input=2.349609375, output=-0.702435103889
			11'd602: out = 32'b10000000000000000101101001000100; // input=2.353515625, output=-0.705210002498
			11'd603: out = 32'b10000000000000000101101010011111; // input=2.357421875, output=-0.707974140471
			11'd604: out = 32'b10000000000000000101101011111001; // input=2.361328125, output=-0.710727475628
			11'd605: out = 32'b10000000000000000101101101010011; // input=2.365234375, output=-0.713469965959
			11'd606: out = 32'b10000000000000000101101110101100; // input=2.369140625, output=-0.716201569616
			11'd607: out = 32'b10000000000000000101110000000110; // input=2.373046875, output=-0.718922244918
			11'd608: out = 32'b10000000000000000101110001011110; // input=2.376953125, output=-0.721631950352
			11'd609: out = 32'b10000000000000000101110010110111; // input=2.380859375, output=-0.724330644569
			11'd610: out = 32'b10000000000000000101110100001111; // input=2.384765625, output=-0.727018286392
			11'd611: out = 32'b10000000000000000101110101100111; // input=2.388671875, output=-0.729694834811
			11'd612: out = 32'b10000000000000000101110110111110; // input=2.392578125, output=-0.732360248984
			11'd613: out = 32'b10000000000000000101111000010101; // input=2.396484375, output=-0.735014488241
			11'd614: out = 32'b10000000000000000101111001101100; // input=2.400390625, output=-0.737657512081
			11'd615: out = 32'b10000000000000000101111011000010; // input=2.404296875, output=-0.740289280175
			11'd616: out = 32'b10000000000000000101111100011000; // input=2.408203125, output=-0.742909752365
			11'd617: out = 32'b10000000000000000101111101101101; // input=2.412109375, output=-0.745518888667
			11'd618: out = 32'b10000000000000000101111111000010; // input=2.416015625, output=-0.748116649267
			11'd619: out = 32'b10000000000000000110000000010111; // input=2.419921875, output=-0.750702994528
			11'd620: out = 32'b10000000000000000110000001101011; // input=2.423828125, output=-0.753277884985
			11'd621: out = 32'b10000000000000000110000010111111; // input=2.427734375, output=-0.755841281348
			11'd622: out = 32'b10000000000000000110000100010011; // input=2.431640625, output=-0.758393144503
			11'd623: out = 32'b10000000000000000110000101100110; // input=2.435546875, output=-0.760933435512
			11'd624: out = 32'b10000000000000000110000110111001; // input=2.439453125, output=-0.763462115613
			11'd625: out = 32'b10000000000000000110001000001100; // input=2.443359375, output=-0.765979146221
			11'd626: out = 32'b10000000000000000110001001011110; // input=2.447265625, output=-0.76848448893
			11'd627: out = 32'b10000000000000000110001010101111; // input=2.451171875, output=-0.770978105511
			11'd628: out = 32'b10000000000000000110001100000001; // input=2.455078125, output=-0.773459957915
			11'd629: out = 32'b10000000000000000110001101010010; // input=2.458984375, output=-0.775930008271
			11'd630: out = 32'b10000000000000000110001110100010; // input=2.462890625, output=-0.77838821889
			11'd631: out = 32'b10000000000000000110001111110010; // input=2.466796875, output=-0.780834552263
			11'd632: out = 32'b10000000000000000110010001000010; // input=2.470703125, output=-0.783268971061
			11'd633: out = 32'b10000000000000000110010010010010; // input=2.474609375, output=-0.785691438138
			11'd634: out = 32'b10000000000000000110010011100001; // input=2.478515625, output=-0.78810191653
			11'd635: out = 32'b10000000000000000110010100101111; // input=2.482421875, output=-0.790500369457
			11'd636: out = 32'b10000000000000000110010101111101; // input=2.486328125, output=-0.792886760321
			11'd637: out = 32'b10000000000000000110010111001011; // input=2.490234375, output=-0.795261052708
			11'd638: out = 32'b10000000000000000110011000011001; // input=2.494140625, output=-0.797623210391
			11'd639: out = 32'b10000000000000000110011001100110; // input=2.498046875, output=-0.799973197324
			11'd640: out = 32'b10000000000000000110011010110010; // input=2.501953125, output=-0.802310977651
			11'd641: out = 32'b10000000000000000110011011111110; // input=2.505859375, output=-0.804636515699
			11'd642: out = 32'b10000000000000000110011101001010; // input=2.509765625, output=-0.806949775984
			11'd643: out = 32'b10000000000000000110011110010110; // input=2.513671875, output=-0.809250723208
			11'd644: out = 32'b10000000000000000110011111100001; // input=2.517578125, output=-0.811539322262
			11'd645: out = 32'b10000000000000000110100000101011; // input=2.521484375, output=-0.813815538224
			11'd646: out = 32'b10000000000000000110100001110101; // input=2.525390625, output=-0.816079336362
			11'd647: out = 32'b10000000000000000110100010111111; // input=2.529296875, output=-0.818330682134
			11'd648: out = 32'b10000000000000000110100100001000; // input=2.533203125, output=-0.820569541186
			11'd649: out = 32'b10000000000000000110100101010001; // input=2.537109375, output=-0.822795879357
			11'd650: out = 32'b10000000000000000110100110011010; // input=2.541015625, output=-0.825009662675
			11'd651: out = 32'b10000000000000000110100111100010; // input=2.544921875, output=-0.82721085736
			11'd652: out = 32'b10000000000000000110101000101010; // input=2.548828125, output=-0.829399429826
			11'd653: out = 32'b10000000000000000110101001110001; // input=2.552734375, output=-0.831575346677
			11'd654: out = 32'b10000000000000000110101010111000; // input=2.556640625, output=-0.833738574711
			11'd655: out = 32'b10000000000000000110101011111110; // input=2.560546875, output=-0.83588908092
			11'd656: out = 32'b10000000000000000110101101000100; // input=2.564453125, output=-0.83802683249
			11'd657: out = 32'b10000000000000000110101110001010; // input=2.568359375, output=-0.840151796802
			11'd658: out = 32'b10000000000000000110101111001111; // input=2.572265625, output=-0.842263941431
			11'd659: out = 32'b10000000000000000110110000010100; // input=2.576171875, output=-0.844363234149
			11'd660: out = 32'b10000000000000000110110001011000; // input=2.580078125, output=-0.846449642922
			11'd661: out = 32'b10000000000000000110110010011100; // input=2.583984375, output=-0.848523135916
			11'd662: out = 32'b10000000000000000110110011100000; // input=2.587890625, output=-0.85058368149
			11'd663: out = 32'b10000000000000000110110100100011; // input=2.591796875, output=-0.852631248204
			11'd664: out = 32'b10000000000000000110110101100110; // input=2.595703125, output=-0.854665804814
			11'd665: out = 32'b10000000000000000110110110101000; // input=2.599609375, output=-0.856687320275
			11'd666: out = 32'b10000000000000000110110111101010; // input=2.603515625, output=-0.858695763742
			11'd667: out = 32'b10000000000000000110111000101011; // input=2.607421875, output=-0.860691104568
			11'd668: out = 32'b10000000000000000110111001101100; // input=2.611328125, output=-0.862673312307
			11'd669: out = 32'b10000000000000000110111010101101; // input=2.615234375, output=-0.864642356712
			11'd670: out = 32'b10000000000000000110111011101101; // input=2.619140625, output=-0.866598207739
			11'd671: out = 32'b10000000000000000110111100101100; // input=2.623046875, output=-0.868540835543
			11'd672: out = 32'b10000000000000000110111101101100; // input=2.626953125, output=-0.870470210483
			11'd673: out = 32'b10000000000000000110111110101010; // input=2.630859375, output=-0.872386303118
			11'd674: out = 32'b10000000000000000110111111101001; // input=2.634765625, output=-0.874289084212
			11'd675: out = 32'b10000000000000000111000000100111; // input=2.638671875, output=-0.87617852473
			11'd676: out = 32'b10000000000000000111000001100100; // input=2.642578125, output=-0.878054595842
			11'd677: out = 32'b10000000000000000111000010100001; // input=2.646484375, output=-0.879917268921
			11'd678: out = 32'b10000000000000000111000011011110; // input=2.650390625, output=-0.881766515544
			11'd679: out = 32'b10000000000000000111000100011010; // input=2.654296875, output=-0.883602307496
			11'd680: out = 32'b10000000000000000111000101010110; // input=2.658203125, output=-0.885424616764
			11'd681: out = 32'b10000000000000000111000110010001; // input=2.662109375, output=-0.887233415541
			11'd682: out = 32'b10000000000000000111000111001100; // input=2.666015625, output=-0.889028676228
			11'd683: out = 32'b10000000000000000111001000000110; // input=2.669921875, output=-0.890810371432
			11'd684: out = 32'b10000000000000000111001001000000; // input=2.673828125, output=-0.892578473965
			11'd685: out = 32'b10000000000000000111001001111010; // input=2.677734375, output=-0.894332956848
			11'd686: out = 32'b10000000000000000111001010110011; // input=2.681640625, output=-0.896073793311
			11'd687: out = 32'b10000000000000000111001011101011; // input=2.685546875, output=-0.897800956791
			11'd688: out = 32'b10000000000000000111001100100011; // input=2.689453125, output=-0.899514420932
			11'd689: out = 32'b10000000000000000111001101011011; // input=2.693359375, output=-0.90121415959
			11'd690: out = 32'b10000000000000000111001110010010; // input=2.697265625, output=-0.902900146829
			11'd691: out = 32'b10000000000000000111001111001001; // input=2.701171875, output=-0.904572356923
			11'd692: out = 32'b10000000000000000111001111111111; // input=2.705078125, output=-0.906230764355
			11'd693: out = 32'b10000000000000000111010000110101; // input=2.708984375, output=-0.907875343821
			11'd694: out = 32'b10000000000000000111010001101011; // input=2.712890625, output=-0.909506070226
			11'd695: out = 32'b10000000000000000111010010100000; // input=2.716796875, output=-0.911122918687
			11'd696: out = 32'b10000000000000000111010011010100; // input=2.720703125, output=-0.912725864533
			11'd697: out = 32'b10000000000000000111010100001000; // input=2.724609375, output=-0.914314883306
			11'd698: out = 32'b10000000000000000111010100111100; // input=2.728515625, output=-0.915889950759
			11'd699: out = 32'b10000000000000000111010101101111; // input=2.732421875, output=-0.917451042858
			11'd700: out = 32'b10000000000000000111010110100010; // input=2.736328125, output=-0.918998135783
			11'd701: out = 32'b10000000000000000111010111010100; // input=2.740234375, output=-0.920531205927
			11'd702: out = 32'b10000000000000000111011000000110; // input=2.744140625, output=-0.922050229897
			11'd703: out = 32'b10000000000000000111011000110111; // input=2.748046875, output=-0.923555184515
			11'd704: out = 32'b10000000000000000111011001101000; // input=2.751953125, output=-0.925046046817
			11'd705: out = 32'b10000000000000000111011010011000; // input=2.755859375, output=-0.926522794055
			11'd706: out = 32'b10000000000000000111011011001000; // input=2.759765625, output=-0.927985403695
			11'd707: out = 32'b10000000000000000111011011111000; // input=2.763671875, output=-0.929433853419
			11'd708: out = 32'b10000000000000000111011100100111; // input=2.767578125, output=-0.930868121127
			11'd709: out = 32'b10000000000000000111011101010101; // input=2.771484375, output=-0.932288184932
			11'd710: out = 32'b10000000000000000111011110000011; // input=2.775390625, output=-0.933694023166
			11'd711: out = 32'b10000000000000000111011110110001; // input=2.779296875, output=-0.935085614378
			11'd712: out = 32'b10000000000000000111011111011110; // input=2.783203125, output=-0.936462937335
			11'd713: out = 32'b10000000000000000111100000001011; // input=2.787109375, output=-0.937825971019
			11'd714: out = 32'b10000000000000000111100000110111; // input=2.791015625, output=-0.939174694632
			11'd715: out = 32'b10000000000000000111100001100011; // input=2.794921875, output=-0.940509087596
			11'd716: out = 32'b10000000000000000111100010001110; // input=2.798828125, output=-0.941829129547
			11'd717: out = 32'b10000000000000000111100010111001; // input=2.802734375, output=-0.943134800345
			11'd718: out = 32'b10000000000000000111100011100011; // input=2.806640625, output=-0.944426080067
			11'd719: out = 32'b10000000000000000111100100001101; // input=2.810546875, output=-0.945702949008
			11'd720: out = 32'b10000000000000000111100100110110; // input=2.814453125, output=-0.946965387686
			11'd721: out = 32'b10000000000000000111100101011111; // input=2.818359375, output=-0.948213376837
			11'd722: out = 32'b10000000000000000111100110000111; // input=2.822265625, output=-0.949446897419
			11'd723: out = 32'b10000000000000000111100110101111; // input=2.826171875, output=-0.950665930609
			11'd724: out = 32'b10000000000000000111100111010111; // input=2.830078125, output=-0.951870457806
			11'd725: out = 32'b10000000000000000111100111111110; // input=2.833984375, output=-0.953060460632
			11'd726: out = 32'b10000000000000000111101000100100; // input=2.837890625, output=-0.954235920927
			11'd727: out = 32'b10000000000000000111101001001010; // input=2.841796875, output=-0.955396820757
			11'd728: out = 32'b10000000000000000111101001110000; // input=2.845703125, output=-0.956543142406
			11'd729: out = 32'b10000000000000000111101010010101; // input=2.849609375, output=-0.957674868384
			11'd730: out = 32'b10000000000000000111101010111010; // input=2.853515625, output=-0.958791981422
			11'd731: out = 32'b10000000000000000111101011011110; // input=2.857421875, output=-0.959894464473
			11'd732: out = 32'b10000000000000000111101100000001; // input=2.861328125, output=-0.960982300717
			11'd733: out = 32'b10000000000000000111101100100101; // input=2.865234375, output=-0.962055473552
			11'd734: out = 32'b10000000000000000111101101000111; // input=2.869140625, output=-0.963113966605
			11'd735: out = 32'b10000000000000000111101101101010; // input=2.873046875, output=-0.964157763723
			11'd736: out = 32'b10000000000000000111101110001011; // input=2.876953125, output=-0.965186848981
			11'd737: out = 32'b10000000000000000111101110101100; // input=2.880859375, output=-0.966201206674
			11'd738: out = 32'b10000000000000000111101111001101; // input=2.884765625, output=-0.967200821326
			11'd739: out = 32'b10000000000000000111101111101110; // input=2.888671875, output=-0.968185677683
			11'd740: out = 32'b10000000000000000111110000001101; // input=2.892578125, output=-0.969155760718
			11'd741: out = 32'b10000000000000000111110000101101; // input=2.896484375, output=-0.970111055629
			11'd742: out = 32'b10000000000000000111110001001011; // input=2.900390625, output=-0.971051547838
			11'd743: out = 32'b10000000000000000111110001101010; // input=2.904296875, output=-0.971977222996
			11'd744: out = 32'b10000000000000000111110010001000; // input=2.908203125, output=-0.972888066977
			11'd745: out = 32'b10000000000000000111110010100101; // input=2.912109375, output=-0.973784065883
			11'd746: out = 32'b10000000000000000111110011000010; // input=2.916015625, output=-0.974665206042
			11'd747: out = 32'b10000000000000000111110011011110; // input=2.919921875, output=-0.975531474009
			11'd748: out = 32'b10000000000000000111110011111010; // input=2.923828125, output=-0.976382856567
			11'd749: out = 32'b10000000000000000111110100010110; // input=2.927734375, output=-0.977219340723
			11'd750: out = 32'b10000000000000000111110100110000; // input=2.931640625, output=-0.978040913714
			11'd751: out = 32'b10000000000000000111110101001011; // input=2.935546875, output=-0.978847563005
			11'd752: out = 32'b10000000000000000111110101100101; // input=2.939453125, output=-0.979639276285
			11'd753: out = 32'b10000000000000000111110101111110; // input=2.943359375, output=-0.980416041476
			11'd754: out = 32'b10000000000000000111110110010111; // input=2.947265625, output=-0.981177846724
			11'd755: out = 32'b10000000000000000111110110110000; // input=2.951171875, output=-0.981924680406
			11'd756: out = 32'b10000000000000000111110111001000; // input=2.955078125, output=-0.982656531125
			11'd757: out = 32'b10000000000000000111110111011111; // input=2.958984375, output=-0.983373387714
			11'd758: out = 32'b10000000000000000111110111110110; // input=2.962890625, output=-0.984075239235
			11'd759: out = 32'b10000000000000000111111000001101; // input=2.966796875, output=-0.984762074979
			11'd760: out = 32'b10000000000000000111111000100011; // input=2.970703125, output=-0.985433884466
			11'd761: out = 32'b10000000000000000111111000111000; // input=2.974609375, output=-0.986090657443
			11'd762: out = 32'b10000000000000000111111001001101; // input=2.978515625, output=-0.986732383891
			11'd763: out = 32'b10000000000000000111111001100010; // input=2.982421875, output=-0.987359054016
			11'd764: out = 32'b10000000000000000111111001110110; // input=2.986328125, output=-0.987970658257
			11'd765: out = 32'b10000000000000000111111010001001; // input=2.990234375, output=-0.988567187281
			11'd766: out = 32'b10000000000000000111111010011100; // input=2.994140625, output=-0.989148631986
			11'd767: out = 32'b10000000000000000111111010101111; // input=2.998046875, output=-0.9897149835
			11'd768: out = 32'b10000000000000000111111011000001; // input=3.001953125, output=-0.990266233181
			11'd769: out = 32'b10000000000000000111111011010011; // input=3.005859375, output=-0.990802372617
			11'd770: out = 32'b10000000000000000111111011100100; // input=3.009765625, output=-0.991323393629
			11'd771: out = 32'b10000000000000000111111011110100; // input=3.013671875, output=-0.991829288265
			11'd772: out = 32'b10000000000000000111111100000100; // input=3.017578125, output=-0.992320048806
			11'd773: out = 32'b10000000000000000111111100010100; // input=3.021484375, output=-0.992795667765
			11'd774: out = 32'b10000000000000000111111100100011; // input=3.025390625, output=-0.993256137883
			11'd775: out = 32'b10000000000000000111111100110010; // input=3.029296875, output=-0.993701452134
			11'd776: out = 32'b10000000000000000111111101000000; // input=3.033203125, output=-0.994131603724
			11'd777: out = 32'b10000000000000000111111101001101; // input=3.037109375, output=-0.994546586089
			11'd778: out = 32'b10000000000000000111111101011010; // input=3.041015625, output=-0.994946392896
			11'd779: out = 32'b10000000000000000111111101100111; // input=3.044921875, output=-0.995331018046
			11'd780: out = 32'b10000000000000000111111101110011; // input=3.048828125, output=-0.995700455669
			11'd781: out = 32'b10000000000000000111111101111111; // input=3.052734375, output=-0.996054700128
			11'd782: out = 32'b10000000000000000111111110001010; // input=3.056640625, output=-0.996393746017
			11'd783: out = 32'b10000000000000000111111110010100; // input=3.060546875, output=-0.996717588164
			11'd784: out = 32'b10000000000000000111111110011111; // input=3.064453125, output=-0.997026221627
			11'd785: out = 32'b10000000000000000111111110101000; // input=3.068359375, output=-0.997319641697
			11'd786: out = 32'b10000000000000000111111110110001; // input=3.072265625, output=-0.997597843896
			11'd787: out = 32'b10000000000000000111111110111010; // input=3.076171875, output=-0.997860823979
			11'd788: out = 32'b10000000000000000111111111000010; // input=3.080078125, output=-0.998108577933
			11'd789: out = 32'b10000000000000000111111111001010; // input=3.083984375, output=-0.998341101979
			11'd790: out = 32'b10000000000000000111111111010001; // input=3.087890625, output=-0.998558392568
			11'd791: out = 32'b10000000000000000111111111010111; // input=3.091796875, output=-0.998760446384
			11'd792: out = 32'b10000000000000000111111111011110; // input=3.095703125, output=-0.998947260345
			11'd793: out = 32'b10000000000000000111111111100011; // input=3.099609375, output=-0.999118831599
			11'd794: out = 32'b10000000000000000111111111101000; // input=3.103515625, output=-0.99927515753
			11'd795: out = 32'b10000000000000000111111111101101; // input=3.107421875, output=-0.999416235751
			11'd796: out = 32'b10000000000000000111111111110001; // input=3.111328125, output=-0.99954206411
			11'd797: out = 32'b10000000000000000111111111110101; // input=3.115234375, output=-0.999652640687
			11'd798: out = 32'b10000000000000000111111111111000; // input=3.119140625, output=-0.999747963794
			11'd799: out = 32'b10000000000000000111111111111010; // input=3.123046875, output=-0.999828031977
			11'd800: out = 32'b10000000000000000111111111111100; // input=3.126953125, output=-0.999892844015
			11'd801: out = 32'b10000000000000000111111111111110; // input=3.130859375, output=-0.999942398918
			11'd802: out = 32'b10000000000000000111111111111111; // input=3.134765625, output=-0.999976695931
			11'd803: out = 32'b10000000000000000111111111111111; // input=3.138671875, output=-0.999995734529
			11'd804: out = 32'b10000000000000000111111111111111; // input=3.142578125, output=-0.999999514423
			11'd805: out = 32'b10000000000000000111111111111111; // input=3.146484375, output=-0.999988035555
			11'd806: out = 32'b10000000000000000111111111111111; // input=3.150390625, output=-0.999961298099
			11'd807: out = 32'b10000000000000000111111111111101; // input=3.154296875, output=-0.999919302465
			11'd808: out = 32'b10000000000000000111111111111011; // input=3.158203125, output=-0.999862049292
			11'd809: out = 32'b10000000000000000111111111111001; // input=3.162109375, output=-0.999789539454
			11'd810: out = 32'b10000000000000000111111111110110; // input=3.166015625, output=-0.999701774058
			11'd811: out = 32'b10000000000000000111111111110011; // input=3.169921875, output=-0.999598754443
			11'd812: out = 32'b10000000000000000111111111101111; // input=3.173828125, output=-0.999480482181
			11'd813: out = 32'b10000000000000000111111111101011; // input=3.177734375, output=-0.999346959076
			11'd814: out = 32'b10000000000000000111111111100110; // input=3.181640625, output=-0.999198187167
			11'd815: out = 32'b10000000000000000111111111100000; // input=3.185546875, output=-0.999034168722
			11'd816: out = 32'b10000000000000000111111111011010; // input=3.189453125, output=-0.998854906245
			11'd817: out = 32'b10000000000000000111111111010100; // input=3.193359375, output=-0.998660402471
			11'd818: out = 32'b10000000000000000111111111001101; // input=3.197265625, output=-0.998450660368
			11'd819: out = 32'b10000000000000000111111111000110; // input=3.201171875, output=-0.998225683137
			11'd820: out = 32'b10000000000000000111111110111110; // input=3.205078125, output=-0.997985474209
			11'd821: out = 32'b10000000000000000111111110110110; // input=3.208984375, output=-0.997730037251
			11'd822: out = 32'b10000000000000000111111110101101; // input=3.212890625, output=-0.997459376161
			11'd823: out = 32'b10000000000000000111111110100011; // input=3.216796875, output=-0.997173495067
			11'd824: out = 32'b10000000000000000111111110011010; // input=3.220703125, output=-0.996872398333
			11'd825: out = 32'b10000000000000000111111110001111; // input=3.224609375, output=-0.996556090553
			11'd826: out = 32'b10000000000000000111111110000100; // input=3.228515625, output=-0.996224576552
			11'd827: out = 32'b10000000000000000111111101111001; // input=3.232421875, output=-0.995877861391
			11'd828: out = 32'b10000000000000000111111101101101; // input=3.236328125, output=-0.995515950358
			11'd829: out = 32'b10000000000000000111111101100001; // input=3.240234375, output=-0.995138848977
			11'd830: out = 32'b10000000000000000111111101010100; // input=3.244140625, output=-0.994746563001
			11'd831: out = 32'b10000000000000000111111101000111; // input=3.248046875, output=-0.994339098417
			11'd832: out = 32'b10000000000000000111111100111001; // input=3.251953125, output=-0.993916461441
			11'd833: out = 32'b10000000000000000111111100101010; // input=3.255859375, output=-0.993478658524
			11'd834: out = 32'b10000000000000000111111100011011; // input=3.259765625, output=-0.993025696344
			11'd835: out = 32'b10000000000000000111111100001100; // input=3.263671875, output=-0.992557581813
			11'd836: out = 32'b10000000000000000111111011111100; // input=3.267578125, output=-0.992074322076
			11'd837: out = 32'b10000000000000000111111011101100; // input=3.271484375, output=-0.991575924504
			11'd838: out = 32'b10000000000000000111111011011011; // input=3.275390625, output=-0.991062396704
			11'd839: out = 32'b10000000000000000111111011001010; // input=3.279296875, output=-0.990533746511
			11'd840: out = 32'b10000000000000000111111010111000; // input=3.283203125, output=-0.989989981992
			11'd841: out = 32'b10000000000000000111111010100110; // input=3.287109375, output=-0.989431111444
			11'd842: out = 32'b10000000000000000111111010010011; // input=3.291015625, output=-0.988857143395
			11'd843: out = 32'b10000000000000000111111010000000; // input=3.294921875, output=-0.988268086602
			11'd844: out = 32'b10000000000000000111111001101100; // input=3.298828125, output=-0.987663950053
			11'd845: out = 32'b10000000000000000111111001010111; // input=3.302734375, output=-0.987044742969
			11'd846: out = 32'b10000000000000000111111001000011; // input=3.306640625, output=-0.986410474795
			11'd847: out = 32'b10000000000000000111111000101101; // input=3.310546875, output=-0.985761155212
			11'd848: out = 32'b10000000000000000111111000011000; // input=3.314453125, output=-0.985096794126
			11'd849: out = 32'b10000000000000000111111000000001; // input=3.318359375, output=-0.984417401675
			11'd850: out = 32'b10000000000000000111110111101011; // input=3.322265625, output=-0.983722988226
			11'd851: out = 32'b10000000000000000111110111010011; // input=3.326171875, output=-0.983013564374
			11'd852: out = 32'b10000000000000000111110110111100; // input=3.330078125, output=-0.982289140945
			11'd853: out = 32'b10000000000000000111110110100011; // input=3.333984375, output=-0.981549728992
			11'd854: out = 32'b10000000000000000111110110001011; // input=3.337890625, output=-0.980795339798
			11'd855: out = 32'b10000000000000000111110101110001; // input=3.341796875, output=-0.980025984873
			11'd856: out = 32'b10000000000000000111110101011000; // input=3.345703125, output=-0.979241675958
			11'd857: out = 32'b10000000000000000111110100111110; // input=3.349609375, output=-0.978442425019
			11'd858: out = 32'b10000000000000000111110100100011; // input=3.353515625, output=-0.977628244254
			11'd859: out = 32'b10000000000000000111110100001000; // input=3.357421875, output=-0.976799146083
			11'd860: out = 32'b10000000000000000111110011101100; // input=3.361328125, output=-0.97595514316
			11'd861: out = 32'b10000000000000000111110011010000; // input=3.365234375, output=-0.975096248362
			11'd862: out = 32'b10000000000000000111110010110011; // input=3.369140625, output=-0.974222474795
			11'd863: out = 32'b10000000000000000111110010010110; // input=3.373046875, output=-0.973333835791
			11'd864: out = 32'b10000000000000000111110001111001; // input=3.376953125, output=-0.972430344911
			11'd865: out = 32'b10000000000000000111110001011011; // input=3.380859375, output=-0.97151201594
			11'd866: out = 32'b10000000000000000111110000111100; // input=3.384765625, output=-0.970578862891
			11'd867: out = 32'b10000000000000000111110000011101; // input=3.388671875, output=-0.969630900003
			11'd868: out = 32'b10000000000000000111101111111101; // input=3.392578125, output=-0.96866814174
			11'd869: out = 32'b10000000000000000111101111011101; // input=3.396484375, output=-0.967690602793
			11'd870: out = 32'b10000000000000000111101110111101; // input=3.400390625, output=-0.966698298078
			11'd871: out = 32'b10000000000000000111101110011100; // input=3.404296875, output=-0.965691242737
			11'd872: out = 32'b10000000000000000111101101111010; // input=3.408203125, output=-0.964669452135
			11'd873: out = 32'b10000000000000000111101101011000; // input=3.412109375, output=-0.963632941864
			11'd874: out = 32'b10000000000000000111101100110110; // input=3.416015625, output=-0.96258172774
			11'd875: out = 32'b10000000000000000111101100010011; // input=3.419921875, output=-0.961515825803
			11'd876: out = 32'b10000000000000000111101011110000; // input=3.423828125, output=-0.960435252318
			11'd877: out = 32'b10000000000000000111101011001100; // input=3.427734375, output=-0.959340023773
			11'd878: out = 32'b10000000000000000111101010100111; // input=3.431640625, output=-0.958230156879
			11'd879: out = 32'b10000000000000000111101010000010; // input=3.435546875, output=-0.957105668571
			11'd880: out = 32'b10000000000000000111101001011101; // input=3.439453125, output=-0.955966576009
			11'd881: out = 32'b10000000000000000111101000110111; // input=3.443359375, output=-0.954812896573
			11'd882: out = 32'b10000000000000000111101000010001; // input=3.447265625, output=-0.953644647867
			11'd883: out = 32'b10000000000000000111100111101010; // input=3.451171875, output=-0.952461847717
			11'd884: out = 32'b10000000000000000111100111000011; // input=3.455078125, output=-0.951264514171
			11'd885: out = 32'b10000000000000000111100110011011; // input=3.458984375, output=-0.950052665499
			11'd886: out = 32'b10000000000000000111100101110011; // input=3.462890625, output=-0.948826320192
			11'd887: out = 32'b10000000000000000111100101001010; // input=3.466796875, output=-0.947585496963
			11'd888: out = 32'b10000000000000000111100100100001; // input=3.470703125, output=-0.946330214745
			11'd889: out = 32'b10000000000000000111100011111000; // input=3.474609375, output=-0.945060492692
			11'd890: out = 32'b10000000000000000111100011001110; // input=3.478515625, output=-0.943776350179
			11'd891: out = 32'b10000000000000000111100010100011; // input=3.482421875, output=-0.9424778068
			11'd892: out = 32'b10000000000000000111100001111000; // input=3.486328125, output=-0.94116488237
			11'd893: out = 32'b10000000000000000111100001001101; // input=3.490234375, output=-0.939837596921
			11'd894: out = 32'b10000000000000000111100000100001; // input=3.494140625, output=-0.938495970706
			11'd895: out = 32'b10000000000000000111011111110100; // input=3.498046875, output=-0.937140024198
			11'd896: out = 32'b10000000000000000111011111000111; // input=3.501953125, output=-0.935769778086
			11'd897: out = 32'b10000000000000000111011110011010; // input=3.505859375, output=-0.934385253279
			11'd898: out = 32'b10000000000000000111011101101100; // input=3.509765625, output=-0.932986470902
			11'd899: out = 32'b10000000000000000111011100111110; // input=3.513671875, output=-0.931573452299
			11'd900: out = 32'b10000000000000000111011100001111; // input=3.517578125, output=-0.930146219032
			11'd901: out = 32'b10000000000000000111011011100000; // input=3.521484375, output=-0.928704792878
			11'd902: out = 32'b10000000000000000111011010110000; // input=3.525390625, output=-0.927249195831
			11'd903: out = 32'b10000000000000000111011010000000; // input=3.529296875, output=-0.925779450103
			11'd904: out = 32'b10000000000000000111011001001111; // input=3.533203125, output=-0.924295578119
			11'd905: out = 32'b10000000000000000111011000011110; // input=3.537109375, output=-0.922797602521
			11'd906: out = 32'b10000000000000000111010111101101; // input=3.541015625, output=-0.921285546168
			11'd907: out = 32'b10000000000000000111010110111011; // input=3.544921875, output=-0.919759432131
			11'd908: out = 32'b10000000000000000111010110001000; // input=3.548828125, output=-0.918219283696
			11'd909: out = 32'b10000000000000000111010101010101; // input=3.552734375, output=-0.916665124365
			11'd910: out = 32'b10000000000000000111010100100010; // input=3.556640625, output=-0.915096977852
			11'd911: out = 32'b10000000000000000111010011101110; // input=3.560546875, output=-0.913514868085
			11'd912: out = 32'b10000000000000000111010010111010; // input=3.564453125, output=-0.911918819205
			11'd913: out = 32'b10000000000000000111010010000101; // input=3.568359375, output=-0.910308855566
			11'd914: out = 32'b10000000000000000111010001010000; // input=3.572265625, output=-0.908685001733
			11'd915: out = 32'b10000000000000000111010000011010; // input=3.576171875, output=-0.907047282486
			11'd916: out = 32'b10000000000000000111001111100100; // input=3.580078125, output=-0.905395722813
			11'd917: out = 32'b10000000000000000111001110101101; // input=3.583984375, output=-0.903730347915
			11'd918: out = 32'b10000000000000000111001101110110; // input=3.587890625, output=-0.902051183204
			11'd919: out = 32'b10000000000000000111001100111111; // input=3.591796875, output=-0.900358254301
			11'd920: out = 32'b10000000000000000111001100000111; // input=3.595703125, output=-0.89865158704
			11'd921: out = 32'b10000000000000000111001011001111; // input=3.599609375, output=-0.896931207461
			11'd922: out = 32'b10000000000000000111001010010110; // input=3.603515625, output=-0.895197141815
			11'd923: out = 32'b10000000000000000111001001011101; // input=3.607421875, output=-0.893449416562
			11'd924: out = 32'b10000000000000000111001000100011; // input=3.611328125, output=-0.89168805837
			11'd925: out = 32'b10000000000000000111000111101001; // input=3.615234375, output=-0.889913094116
			11'd926: out = 32'b10000000000000000111000110101110; // input=3.619140625, output=-0.888124550883
			11'd927: out = 32'b10000000000000000111000101110011; // input=3.623046875, output=-0.886322455962
			11'd928: out = 32'b10000000000000000111000100111000; // input=3.626953125, output=-0.88450683685
			11'd929: out = 32'b10000000000000000111000011111100; // input=3.630859375, output=-0.882677721253
			11'd930: out = 32'b10000000000000000111000010111111; // input=3.634765625, output=-0.880835137079
			11'd931: out = 32'b10000000000000000111000010000010; // input=3.638671875, output=-0.878979112445
			11'd932: out = 32'b10000000000000000111000001000101; // input=3.642578125, output=-0.877109675671
			11'd933: out = 32'b10000000000000000111000000000111; // input=3.646484375, output=-0.875226855283
			11'd934: out = 32'b10000000000000000110111111001001; // input=3.650390625, output=-0.87333068001
			11'd935: out = 32'b10000000000000000110111110001011; // input=3.654296875, output=-0.871421178785
			11'd936: out = 32'b10000000000000000110111101001100; // input=3.658203125, output=-0.869498380745
			11'd937: out = 32'b10000000000000000110111100001100; // input=3.662109375, output=-0.867562315229
			11'd938: out = 32'b10000000000000000110111011001100; // input=3.666015625, output=-0.86561301178
			11'd939: out = 32'b10000000000000000110111010001100; // input=3.669921875, output=-0.863650500142
			11'd940: out = 32'b10000000000000000110111001001011; // input=3.673828125, output=-0.861674810259
			11'd941: out = 32'b10000000000000000110111000001010; // input=3.677734375, output=-0.859685972279
			11'd942: out = 32'b10000000000000000110110111001001; // input=3.681640625, output=-0.857684016548
			11'd943: out = 32'b10000000000000000110110110000111; // input=3.685546875, output=-0.855668973615
			11'd944: out = 32'b10000000000000000110110101000100; // input=3.689453125, output=-0.853640874226
			11'd945: out = 32'b10000000000000000110110100000001; // input=3.693359375, output=-0.851599749328
			11'd946: out = 32'b10000000000000000110110010111110; // input=3.697265625, output=-0.849545630065
			11'd947: out = 32'b10000000000000000110110001111010; // input=3.701171875, output=-0.847478547781
			11'd948: out = 32'b10000000000000000110110000110110; // input=3.705078125, output=-0.845398534017
			11'd949: out = 32'b10000000000000000110101111110001; // input=3.708984375, output=-0.843305620512
			11'd950: out = 32'b10000000000000000110101110101100; // input=3.712890625, output=-0.8411998392
			11'd951: out = 32'b10000000000000000110101101100111; // input=3.716796875, output=-0.839081222214
			11'd952: out = 32'b10000000000000000110101100100001; // input=3.720703125, output=-0.83694980188
			11'd953: out = 32'b10000000000000000110101011011011; // input=3.724609375, output=-0.834805610723
			11'd954: out = 32'b10000000000000000110101010010100; // input=3.728515625, output=-0.832648681459
			11'd955: out = 32'b10000000000000000110101001001101; // input=3.732421875, output=-0.830479047
			11'd956: out = 32'b10000000000000000110101000000110; // input=3.736328125, output=-0.828296740453
			11'd957: out = 32'b10000000000000000110100110111110; // input=3.740234375, output=-0.826101795117
			11'd958: out = 32'b10000000000000000110100101110101; // input=3.744140625, output=-0.823894244484
			11'd959: out = 32'b10000000000000000110100100101101; // input=3.748046875, output=-0.821674122238
			11'd960: out = 32'b10000000000000000110100011100011; // input=3.751953125, output=-0.819441462256
			11'd961: out = 32'b10000000000000000110100010011010; // input=3.755859375, output=-0.817196298606
			11'd962: out = 32'b10000000000000000110100001010000; // input=3.759765625, output=-0.814938665546
			11'd963: out = 32'b10000000000000000110100000000110; // input=3.763671875, output=-0.812668597524
			11'd964: out = 32'b10000000000000000110011110111011; // input=3.767578125, output=-0.810386129179
			11'd965: out = 32'b10000000000000000110011101110000; // input=3.771484375, output=-0.808091295339
			11'd966: out = 32'b10000000000000000110011100100100; // input=3.775390625, output=-0.80578413102
			11'd967: out = 32'b10000000000000000110011011011000; // input=3.779296875, output=-0.803464671426
			11'd968: out = 32'b10000000000000000110011010001100; // input=3.783203125, output=-0.801132951951
			11'd969: out = 32'b10000000000000000110011000111111; // input=3.787109375, output=-0.798789008172
			11'd970: out = 32'b10000000000000000110010111110010; // input=3.791015625, output=-0.796432875855
			11'd971: out = 32'b10000000000000000110010110100100; // input=3.794921875, output=-0.794064590953
			11'd972: out = 32'b10000000000000000110010101010110; // input=3.798828125, output=-0.791684189602
			11'd973: out = 32'b10000000000000000110010100001000; // input=3.802734375, output=-0.789291708124
			11'd974: out = 32'b10000000000000000110010010111001; // input=3.806640625, output=-0.786887183026
			11'd975: out = 32'b10000000000000000110010001101010; // input=3.810546875, output=-0.784470650998
			11'd976: out = 32'b10000000000000000110010000011010; // input=3.814453125, output=-0.782042148913
			11'd977: out = 32'b10000000000000000110001111001010; // input=3.818359375, output=-0.779601713826
			11'd978: out = 32'b10000000000000000110001101111010; // input=3.822265625, output=-0.777149382977
			11'd979: out = 32'b10000000000000000110001100101001; // input=3.826171875, output=-0.774685193784
			11'd980: out = 32'b10000000000000000110001011011000; // input=3.830078125, output=-0.772209183849
			11'd981: out = 32'b10000000000000000110001010000110; // input=3.833984375, output=-0.769721390951
			11'd982: out = 32'b10000000000000000110001000110100; // input=3.837890625, output=-0.767221853052
			11'd983: out = 32'b10000000000000000110000111100010; // input=3.841796875, output=-0.764710608291
			11'd984: out = 32'b10000000000000000110000110001111; // input=3.845703125, output=-0.762187694988
			11'd985: out = 32'b10000000000000000110000100111100; // input=3.849609375, output=-0.759653151638
			11'd986: out = 32'b10000000000000000110000011101001; // input=3.853515625, output=-0.757107016915
			11'd987: out = 32'b10000000000000000110000010010101; // input=3.857421875, output=-0.754549329671
			11'd988: out = 32'b10000000000000000110000001000001; // input=3.861328125, output=-0.751980128932
			11'd989: out = 32'b10000000000000000101111111101100; // input=3.865234375, output=-0.749399453902
			11'd990: out = 32'b10000000000000000101111110010111; // input=3.869140625, output=-0.746807343958
			11'd991: out = 32'b10000000000000000101111101000010; // input=3.873046875, output=-0.744203838653
			11'd992: out = 32'b10000000000000000101111011101100; // input=3.876953125, output=-0.741588977713
			11'd993: out = 32'b10000000000000000101111010010110; // input=3.880859375, output=-0.738962801038
			11'd994: out = 32'b10000000000000000101111001000000; // input=3.884765625, output=-0.736325348699
			11'd995: out = 32'b10000000000000000101110111101001; // input=3.888671875, output=-0.733676660942
			11'd996: out = 32'b10000000000000000101110110010010; // input=3.892578125, output=-0.731016778181
			11'd997: out = 32'b10000000000000000101110100111010; // input=3.896484375, output=-0.728345741004
			11'd998: out = 32'b10000000000000000101110011100011; // input=3.900390625, output=-0.725663590167
			11'd999: out = 32'b10000000000000000101110010001010; // input=3.904296875, output=-0.722970366596
			11'd1000: out = 32'b10000000000000000101110000110010; // input=3.908203125, output=-0.720266111387
			11'd1001: out = 32'b10000000000000000101101111011001; // input=3.912109375, output=-0.717550865803
			11'd1002: out = 32'b10000000000000000101101101111111; // input=3.916015625, output=-0.714824671276
			11'd1003: out = 32'b10000000000000000101101100100110; // input=3.919921875, output=-0.712087569404
			11'd1004: out = 32'b10000000000000000101101011001100; // input=3.923828125, output=-0.709339601952
			11'd1005: out = 32'b10000000000000000101101001110001; // input=3.927734375, output=-0.70658081085
			11'd1006: out = 32'b10000000000000000101101000010110; // input=3.931640625, output=-0.703811238194
			11'd1007: out = 32'b10000000000000000101100110111011; // input=3.935546875, output=-0.701030926245
			11'd1008: out = 32'b10000000000000000101100101100000; // input=3.939453125, output=-0.698239917426
			11'd1009: out = 32'b10000000000000000101100100000100; // input=3.943359375, output=-0.695438254325
			11'd1010: out = 32'b10000000000000000101100010101000; // input=3.947265625, output=-0.692625979692
			11'd1011: out = 32'b10000000000000000101100001001011; // input=3.951171875, output=-0.689803136439
			11'd1012: out = 32'b10000000000000000101011111101111; // input=3.955078125, output=-0.686969767639
			11'd1013: out = 32'b10000000000000000101011110010001; // input=3.958984375, output=-0.684125916525
			11'd1014: out = 32'b10000000000000000101011100110100; // input=3.962890625, output=-0.681271626491
			11'd1015: out = 32'b10000000000000000101011011010110; // input=3.966796875, output=-0.678406941091
			11'd1016: out = 32'b10000000000000000101011001111000; // input=3.970703125, output=-0.675531904035
			11'd1017: out = 32'b10000000000000000101011000011001; // input=3.974609375, output=-0.672646559194
			11'd1018: out = 32'b10000000000000000101010110111010; // input=3.978515625, output=-0.669750950593
			11'd1019: out = 32'b10000000000000000101010101011011; // input=3.982421875, output=-0.666845122418
			11'd1020: out = 32'b10000000000000000101010011111100; // input=3.986328125, output=-0.663929119006
			11'd1021: out = 32'b10000000000000000101010010011100; // input=3.990234375, output=-0.661002984852
			11'd1022: out = 32'b10000000000000000101010000111100; // input=3.994140625, output=-0.658066764607
			11'd1023: out = 32'b10000000000000000101001111011011; // input=3.998046875, output=-0.655120503072
			11'd1024: out = 32'b00000000000000000111111111111111; // input=-0.001953125, output=0.999998092652
			11'd1025: out = 32'b00000000000000000111111111111111; // input=-0.005859375, output=0.999982833911
			11'd1026: out = 32'b00000000000000000111111111111110; // input=-0.009765625, output=0.999952316663
			11'd1027: out = 32'b00000000000000000111111111111101; // input=-0.013671875, output=0.999906541373
			11'd1028: out = 32'b00000000000000000111111111111011; // input=-0.017578125, output=0.999845508739
			11'd1029: out = 32'b00000000000000000111111111111000; // input=-0.021484375, output=0.999769219693
			11'd1030: out = 32'b00000000000000000111111111110101; // input=-0.025390625, output=0.999677675398
			11'd1031: out = 32'b00000000000000000111111111110010; // input=-0.029296875, output=0.999570877252
			11'd1032: out = 32'b00000000000000000111111111101110; // input=-0.033203125, output=0.999448826885
			11'd1033: out = 32'b00000000000000000111111111101001; // input=-0.037109375, output=0.999311526157
			11'd1034: out = 32'b00000000000000000111111111100100; // input=-0.041015625, output=0.999158977166
			11'd1035: out = 32'b00000000000000000111111111011111; // input=-0.044921875, output=0.998991182238
			11'd1036: out = 32'b00000000000000000111111111011001; // input=-0.048828125, output=0.998808143933
			11'd1037: out = 32'b00000000000000000111111111010010; // input=-0.052734375, output=0.998609865045
			11'd1038: out = 32'b00000000000000000111111111001011; // input=-0.056640625, output=0.998396348599
			11'd1039: out = 32'b00000000000000000111111111000100; // input=-0.060546875, output=0.998167597854
			11'd1040: out = 32'b00000000000000000111111110111100; // input=-0.064453125, output=0.997923616299
			11'd1041: out = 32'b00000000000000000111111110110011; // input=-0.068359375, output=0.997664407657
			11'd1042: out = 32'b00000000000000000111111110101010; // input=-0.072265625, output=0.997389975884
			11'd1043: out = 32'b00000000000000000111111110100001; // input=-0.076171875, output=0.997100325166
			11'd1044: out = 32'b00000000000000000111111110010111; // input=-0.080078125, output=0.996795459925
			11'd1045: out = 32'b00000000000000000111111110001101; // input=-0.083984375, output=0.996475384812
			11'd1046: out = 32'b00000000000000000111111110000010; // input=-0.087890625, output=0.99614010471
			11'd1047: out = 32'b00000000000000000111111101110110; // input=-0.091796875, output=0.995789624735
			11'd1048: out = 32'b00000000000000000111111101101010; // input=-0.095703125, output=0.995423950236
			11'd1049: out = 32'b00000000000000000111111101011110; // input=-0.099609375, output=0.995043086793
			11'd1050: out = 32'b00000000000000000111111101010001; // input=-0.103515625, output=0.994647040216
			11'd1051: out = 32'b00000000000000000111111101000011; // input=-0.107421875, output=0.994235816549
			11'd1052: out = 32'b00000000000000000111111100110101; // input=-0.111328125, output=0.993809422066
			11'd1053: out = 32'b00000000000000000111111100100111; // input=-0.115234375, output=0.993367863275
			11'd1054: out = 32'b00000000000000000111111100011000; // input=-0.119140625, output=0.992911146912
			11'd1055: out = 32'b00000000000000000111111100001000; // input=-0.123046875, output=0.992439279947
			11'd1056: out = 32'b00000000000000000111111011111000; // input=-0.126953125, output=0.991952269579
			11'd1057: out = 32'b00000000000000000111111011101000; // input=-0.130859375, output=0.99145012324
			11'd1058: out = 32'b00000000000000000111111011010111; // input=-0.134765625, output=0.990932848592
			11'd1059: out = 32'b00000000000000000111111011000101; // input=-0.138671875, output=0.990400453528
			11'd1060: out = 32'b00000000000000000111111010110100; // input=-0.142578125, output=0.989852946172
			11'd1061: out = 32'b00000000000000000111111010100001; // input=-0.146484375, output=0.989290334878
			11'd1062: out = 32'b00000000000000000111111010001110; // input=-0.150390625, output=0.98871262823
			11'd1063: out = 32'b00000000000000000111111001111011; // input=-0.154296875, output=0.988119835044
			11'd1064: out = 32'b00000000000000000111111001100111; // input=-0.158203125, output=0.987511964365
			11'd1065: out = 32'b00000000000000000111111001010010; // input=-0.162109375, output=0.986889025468
			11'd1066: out = 32'b00000000000000000111111000111101; // input=-0.166015625, output=0.986251027859
			11'd1067: out = 32'b00000000000000000111111000101000; // input=-0.169921875, output=0.985597981273
			11'd1068: out = 32'b00000000000000000111111000010010; // input=-0.173828125, output=0.984929895674
			11'd1069: out = 32'b00000000000000000111110111111100; // input=-0.177734375, output=0.984246781257
			11'd1070: out = 32'b00000000000000000111110111100101; // input=-0.181640625, output=0.983548648445
			11'd1071: out = 32'b00000000000000000111110111001110; // input=-0.185546875, output=0.98283550789
			11'd1072: out = 32'b00000000000000000111110110110110; // input=-0.189453125, output=0.982107370475
			11'd1073: out = 32'b00000000000000000111110110011101; // input=-0.193359375, output=0.98136424731
			11'd1074: out = 32'b00000000000000000111110110000101; // input=-0.197265625, output=0.980606149734
			11'd1075: out = 32'b00000000000000000111110101101011; // input=-0.201171875, output=0.979833089314
			11'd1076: out = 32'b00000000000000000111110101010001; // input=-0.205078125, output=0.979045077847
			11'd1077: out = 32'b00000000000000000111110100110111; // input=-0.208984375, output=0.978242127357
			11'd1078: out = 32'b00000000000000000111110100011100; // input=-0.212890625, output=0.977424250095
			11'd1079: out = 32'b00000000000000000111110100000001; // input=-0.216796875, output=0.976591458542
			11'd1080: out = 32'b00000000000000000111110011100101; // input=-0.220703125, output=0.975743765405
			11'd1081: out = 32'b00000000000000000111110011001001; // input=-0.224609375, output=0.974881183619
			11'd1082: out = 32'b00000000000000000111110010101100; // input=-0.228515625, output=0.974003726345
			11'd1083: out = 32'b00000000000000000111110010001111; // input=-0.232421875, output=0.973111406972
			11'd1084: out = 32'b00000000000000000111110001110001; // input=-0.236328125, output=0.972204239117
			11'd1085: out = 32'b00000000000000000111110001010011; // input=-0.240234375, output=0.971282236621
			11'd1086: out = 32'b00000000000000000111110000110100; // input=-0.244140625, output=0.970345413553
			11'd1087: out = 32'b00000000000000000111110000010101; // input=-0.248046875, output=0.969393784208
			11'd1088: out = 32'b00000000000000000111101111110101; // input=-0.251953125, output=0.968427363107
			11'd1089: out = 32'b00000000000000000111101111010101; // input=-0.255859375, output=0.967446164995
			11'd1090: out = 32'b00000000000000000111101110110101; // input=-0.259765625, output=0.966450204846
			11'd1091: out = 32'b00000000000000000111101110010100; // input=-0.263671875, output=0.965439497855
			11'd1092: out = 32'b00000000000000000111101101110010; // input=-0.267578125, output=0.964414059445
			11'd1093: out = 32'b00000000000000000111101101010000; // input=-0.271484375, output=0.963373905264
			11'd1094: out = 32'b00000000000000000111101100101101; // input=-0.275390625, output=0.962319051181
			11'd1095: out = 32'b00000000000000000111101100001010; // input=-0.279296875, output=0.961249513295
			11'd1096: out = 32'b00000000000000000111101011100111; // input=-0.283203125, output=0.960165307923
			11'd1097: out = 32'b00000000000000000111101011000011; // input=-0.287109375, output=0.95906645161
			11'd1098: out = 32'b00000000000000000111101010011110; // input=-0.291015625, output=0.957952961123
			11'd1099: out = 32'b00000000000000000111101001111001; // input=-0.294921875, output=0.956824853452
			11'd1100: out = 32'b00000000000000000111101001010100; // input=-0.298828125, output=0.955682145811
			11'd1101: out = 32'b00000000000000000111101000101110; // input=-0.302734375, output=0.954524855637
			11'd1102: out = 32'b00000000000000000111101000000111; // input=-0.306640625, output=0.953353000587
			11'd1103: out = 32'b00000000000000000111100111100001; // input=-0.310546875, output=0.952166598544
			11'd1104: out = 32'b00000000000000000111100110111001; // input=-0.314453125, output=0.95096566761
			11'd1105: out = 32'b00000000000000000111100110010001; // input=-0.318359375, output=0.94975022611
			11'd1106: out = 32'b00000000000000000111100101101001; // input=-0.322265625, output=0.94852029259
			11'd1107: out = 32'b00000000000000000111100101000000; // input=-0.326171875, output=0.947275885817
			11'd1108: out = 32'b00000000000000000111100100010111; // input=-0.330078125, output=0.94601702478
			11'd1109: out = 32'b00000000000000000111100011101101; // input=-0.333984375, output=0.944743728687
			11'd1110: out = 32'b00000000000000000111100011000011; // input=-0.337890625, output=0.943456016966
			11'd1111: out = 32'b00000000000000000111100010011000; // input=-0.341796875, output=0.942153909268
			11'd1112: out = 32'b00000000000000000111100001101101; // input=-0.345703125, output=0.940837425461
			11'd1113: out = 32'b00000000000000000111100001000010; // input=-0.349609375, output=0.939506585632
			11'd1114: out = 32'b00000000000000000111100000010110; // input=-0.353515625, output=0.938161410088
			11'd1115: out = 32'b00000000000000000111011111101001; // input=-0.357421875, output=0.936801919355
			11'd1116: out = 32'b00000000000000000111011110111100; // input=-0.361328125, output=0.935428134178
			11'd1117: out = 32'b00000000000000000111011110001111; // input=-0.365234375, output=0.934040075518
			11'd1118: out = 32'b00000000000000000111011101100001; // input=-0.369140625, output=0.932637764556
			11'd1119: out = 32'b00000000000000000111011100110010; // input=-0.373046875, output=0.931221222689
			11'd1120: out = 32'b00000000000000000111011100000011; // input=-0.376953125, output=0.929790471532
			11'd1121: out = 32'b00000000000000000111011011010100; // input=-0.380859375, output=0.928345532916
			11'd1122: out = 32'b00000000000000000111011010100100; // input=-0.384765625, output=0.92688642889
			11'd1123: out = 32'b00000000000000000111011001110100; // input=-0.388671875, output=0.925413181717
			11'd1124: out = 32'b00000000000000000111011001000011; // input=-0.392578125, output=0.923925813877
			11'd1125: out = 32'b00000000000000000111011000010010; // input=-0.396484375, output=0.922424348067
			11'd1126: out = 32'b00000000000000000111010111100000; // input=-0.400390625, output=0.920908807195
			11'd1127: out = 32'b00000000000000000111010110101110; // input=-0.404296875, output=0.919379214389
			11'd1128: out = 32'b00000000000000000111010101111100; // input=-0.408203125, output=0.917835592986
			11'd1129: out = 32'b00000000000000000111010101001001; // input=-0.412109375, output=0.916277966542
			11'd1130: out = 32'b00000000000000000111010100010101; // input=-0.416015625, output=0.914706358823
			11'd1131: out = 32'b00000000000000000111010011100001; // input=-0.419921875, output=0.913120793811
			11'd1132: out = 32'b00000000000000000111010010101101; // input=-0.423828125, output=0.911521295699
			11'd1133: out = 32'b00000000000000000111010001111000; // input=-0.427734375, output=0.909907888893
			11'd1134: out = 32'b00000000000000000111010001000011; // input=-0.431640625, output=0.908280598013
			11'd1135: out = 32'b00000000000000000111010000001101; // input=-0.435546875, output=0.906639447888
			11'd1136: out = 32'b00000000000000000111001111010111; // input=-0.439453125, output=0.90498446356
			11'd1137: out = 32'b00000000000000000111001110100000; // input=-0.443359375, output=0.903315670283
			11'd1138: out = 32'b00000000000000000111001101101001; // input=-0.447265625, output=0.901633093521
			11'd1139: out = 32'b00000000000000000111001100110001; // input=-0.451171875, output=0.899936758946
			11'd1140: out = 32'b00000000000000000111001011111001; // input=-0.455078125, output=0.898226692444
			11'd1141: out = 32'b00000000000000000111001011000001; // input=-0.458984375, output=0.896502920108
			11'd1142: out = 32'b00000000000000000111001010001000; // input=-0.462890625, output=0.89476546824
			11'd1143: out = 32'b00000000000000000111001001001110; // input=-0.466796875, output=0.893014363352
			11'd1144: out = 32'b00000000000000000111001000010100; // input=-0.470703125, output=0.891249632163
			11'd1145: out = 32'b00000000000000000111000111011010; // input=-0.474609375, output=0.889471301602
			11'd1146: out = 32'b00000000000000000111000110011111; // input=-0.478515625, output=0.887679398803
			11'd1147: out = 32'b00000000000000000111000101100100; // input=-0.482421875, output=0.885873951108
			11'd1148: out = 32'b00000000000000000111000100101001; // input=-0.486328125, output=0.884054986067
			11'd1149: out = 32'b00000000000000000111000011101101; // input=-0.490234375, output=0.882222531435
			11'd1150: out = 32'b00000000000000000111000010110000; // input=-0.494140625, output=0.880376615172
			11'd1151: out = 32'b00000000000000000111000001110011; // input=-0.498046875, output=0.878517265445
			11'd1152: out = 32'b00000000000000000111000000110110; // input=-0.501953125, output=0.876644510625
			11'd1153: out = 32'b00000000000000000110111111111000; // input=-0.505859375, output=0.874758379289
			11'd1154: out = 32'b00000000000000000110111110111010; // input=-0.509765625, output=0.872858900216
			11'd1155: out = 32'b00000000000000000110111101111011; // input=-0.513671875, output=0.870946102391
			11'd1156: out = 32'b00000000000000000110111100111100; // input=-0.517578125, output=0.869020014999
			11'd1157: out = 32'b00000000000000000110111011111100; // input=-0.521484375, output=0.867080667431
			11'd1158: out = 32'b00000000000000000110111010111101; // input=-0.525390625, output=0.865128089279
			11'd1159: out = 32'b00000000000000000110111001111100; // input=-0.529296875, output=0.863162310337
			11'd1160: out = 32'b00000000000000000110111000111011; // input=-0.533203125, output=0.861183360599
			11'd1161: out = 32'b00000000000000000110110111111010; // input=-0.537109375, output=0.859191270264
			11'd1162: out = 32'b00000000000000000110110110111000; // input=-0.541015625, output=0.857186069726
			11'd1163: out = 32'b00000000000000000110110101110110; // input=-0.544921875, output=0.855167789584
			11'd1164: out = 32'b00000000000000000110110100110100; // input=-0.548828125, output=0.853136460634
			11'd1165: out = 32'b00000000000000000110110011110001; // input=-0.552734375, output=0.85109211387
			11'd1166: out = 32'b00000000000000000110110010101101; // input=-0.556640625, output=0.849034780489
			11'd1167: out = 32'b00000000000000000110110001101001; // input=-0.560546875, output=0.846964491881
			11'd1168: out = 32'b00000000000000000110110000100101; // input=-0.564453125, output=0.844881279637
			11'd1169: out = 32'b00000000000000000110101111100000; // input=-0.568359375, output=0.842785175544
			11'd1170: out = 32'b00000000000000000110101110011011; // input=-0.572265625, output=0.840676211586
			11'd1171: out = 32'b00000000000000000110101101010110; // input=-0.576171875, output=0.838554419944
			11'd1172: out = 32'b00000000000000000110101100010000; // input=-0.580078125, output=0.836419832992
			11'd1173: out = 32'b00000000000000000110101011001001; // input=-0.583984375, output=0.834272483304
			11'd1174: out = 32'b00000000000000000110101010000011; // input=-0.587890625, output=0.832112403643
			11'd1175: out = 32'b00000000000000000110101000111011; // input=-0.591796875, output=0.829939626972
			11'd1176: out = 32'b00000000000000000110100111110100; // input=-0.595703125, output=0.827754186442
			11'd1177: out = 32'b00000000000000000110100110101100; // input=-0.599609375, output=0.825556115402
			11'd1178: out = 32'b00000000000000000110100101100011; // input=-0.603515625, output=0.823345447392
			11'd1179: out = 32'b00000000000000000110100100011011; // input=-0.607421875, output=0.821122216143
			11'd1180: out = 32'b00000000000000000110100011010001; // input=-0.611328125, output=0.818886455579
			11'd1181: out = 32'b00000000000000000110100010001000; // input=-0.615234375, output=0.816638199815
			11'd1182: out = 32'b00000000000000000110100000111110; // input=-0.619140625, output=0.814377483157
			11'd1183: out = 32'b00000000000000000110011111110011; // input=-0.623046875, output=0.812104340101
			11'd1184: out = 32'b00000000000000000110011110101000; // input=-0.626953125, output=0.809818805332
			11'd1185: out = 32'b00000000000000000110011101011101; // input=-0.630859375, output=0.807520913724
			11'd1186: out = 32'b00000000000000000110011100010001; // input=-0.634765625, output=0.80521070034
			11'd1187: out = 32'b00000000000000000110011011000101; // input=-0.638671875, output=0.802888200432
			11'd1188: out = 32'b00000000000000000110011001111001; // input=-0.642578125, output=0.800553449438
			11'd1189: out = 32'b00000000000000000110011000101100; // input=-0.646484375, output=0.798206482983
			11'd1190: out = 32'b00000000000000000110010111011110; // input=-0.650390625, output=0.795847336879
			11'd1191: out = 32'b00000000000000000110010110010001; // input=-0.654296875, output=0.793476047124
			11'd1192: out = 32'b00000000000000000110010101000011; // input=-0.658203125, output=0.791092649901
			11'd1193: out = 32'b00000000000000000110010011110100; // input=-0.662109375, output=0.788697181577
			11'd1194: out = 32'b00000000000000000110010010100101; // input=-0.666015625, output=0.786289678704
			11'd1195: out = 32'b00000000000000000110010001010110; // input=-0.669921875, output=0.783870178019
			11'd1196: out = 32'b00000000000000000110010000000110; // input=-0.673828125, output=0.781438716439
			11'd1197: out = 32'b00000000000000000110001110110110; // input=-0.677734375, output=0.778995331066
			11'd1198: out = 32'b00000000000000000110001101100110; // input=-0.681640625, output=0.776540059182
			11'd1199: out = 32'b00000000000000000110001100010101; // input=-0.685546875, output=0.774072938252
			11'd1200: out = 32'b00000000000000000110001011000100; // input=-0.689453125, output=0.771594005922
			11'd1201: out = 32'b00000000000000000110001001110010; // input=-0.693359375, output=0.769103300017
			11'd1202: out = 32'b00000000000000000110001000100000; // input=-0.697265625, output=0.766600858541
			11'd1203: out = 32'b00000000000000000110000111001110; // input=-0.701171875, output=0.76408671968
			11'd1204: out = 32'b00000000000000000110000101111011; // input=-0.705078125, output=0.761560921795
			11'd1205: out = 32'b00000000000000000110000100101000; // input=-0.708984375, output=0.759023503428
			11'd1206: out = 32'b00000000000000000110000011010100; // input=-0.712890625, output=0.756474503295
			11'd1207: out = 32'b00000000000000000110000010000000; // input=-0.716796875, output=0.753913960293
			11'd1208: out = 32'b00000000000000000110000000101100; // input=-0.720703125, output=0.751341913491
			11'd1209: out = 32'b00000000000000000101111111010111; // input=-0.724609375, output=0.748758402136
			11'd1210: out = 32'b00000000000000000101111110000010; // input=-0.728515625, output=0.746163465649
			11'd1211: out = 32'b00000000000000000101111100101101; // input=-0.732421875, output=0.743557143625
			11'd1212: out = 32'b00000000000000000101111011010111; // input=-0.736328125, output=0.740939475835
			11'd1213: out = 32'b00000000000000000101111010000001; // input=-0.740234375, output=0.738310502219
			11'd1214: out = 32'b00000000000000000101111000101010; // input=-0.744140625, output=0.735670262894
			11'd1215: out = 32'b00000000000000000101110111010100; // input=-0.748046875, output=0.733018798145
			11'd1216: out = 32'b00000000000000000101110101111100; // input=-0.751953125, output=0.730356148432
			11'd1217: out = 32'b00000000000000000101110100100101; // input=-0.755859375, output=0.727682354382
			11'd1218: out = 32'b00000000000000000101110011001101; // input=-0.759765625, output=0.724997456795
			11'd1219: out = 32'b00000000000000000101110001110100; // input=-0.763671875, output=0.722301496639
			11'd1220: out = 32'b00000000000000000101110000011100; // input=-0.767578125, output=0.71959451505
			11'd1221: out = 32'b00000000000000000101101111000011; // input=-0.771484375, output=0.716876553335
			11'd1222: out = 32'b00000000000000000101101101101001; // input=-0.775390625, output=0.714147652965
			11'd1223: out = 32'b00000000000000000101101100001111; // input=-0.779296875, output=0.711407855581
			11'd1224: out = 32'b00000000000000000101101010110101; // input=-0.783203125, output=0.708657202988
			11'd1225: out = 32'b00000000000000000101101001011011; // input=-0.787109375, output=0.705895737158
			11'd1226: out = 32'b00000000000000000101101000000000; // input=-0.791015625, output=0.703123500228
			11'd1227: out = 32'b00000000000000000101100110100101; // input=-0.794921875, output=0.700340534498
			11'd1228: out = 32'b00000000000000000101100101001001; // input=-0.798828125, output=0.697546882433
			11'd1229: out = 32'b00000000000000000101100011101101; // input=-0.802734375, output=0.694742586661
			11'd1230: out = 32'b00000000000000000101100010010001; // input=-0.806640625, output=0.691927689972
			11'd1231: out = 32'b00000000000000000101100000110101; // input=-0.810546875, output=0.689102235318
			11'd1232: out = 32'b00000000000000000101011111011000; // input=-0.814453125, output=0.686266265812
			11'd1233: out = 32'b00000000000000000101011101111010; // input=-0.818359375, output=0.683419824726
			11'd1234: out = 32'b00000000000000000101011100011101; // input=-0.822265625, output=0.680562955495
			11'd1235: out = 32'b00000000000000000101011010111111; // input=-0.826171875, output=0.677695701711
			11'd1236: out = 32'b00000000000000000101011001100000; // input=-0.830078125, output=0.674818107123
			11'd1237: out = 32'b00000000000000000101011000000010; // input=-0.833984375, output=0.671930215642
			11'd1238: out = 32'b00000000000000000101010110100011; // input=-0.837890625, output=0.669032071333
			11'd1239: out = 32'b00000000000000000101010101000100; // input=-0.841796875, output=0.666123718417
			11'd1240: out = 32'b00000000000000000101010011100100; // input=-0.845703125, output=0.663205201273
			11'd1241: out = 32'b00000000000000000101010010000100; // input=-0.849609375, output=0.660276564433
			11'd1242: out = 32'b00000000000000000101010000100100; // input=-0.853515625, output=0.657337852585
			11'd1243: out = 32'b00000000000000000101001111000011; // input=-0.857421875, output=0.654389110571
			11'd1244: out = 32'b00000000000000000101001101100010; // input=-0.861328125, output=0.651430383384
			11'd1245: out = 32'b00000000000000000101001100000001; // input=-0.865234375, output=0.64846171617
			11'd1246: out = 32'b00000000000000000101001010011111; // input=-0.869140625, output=0.645483154229
			11'd1247: out = 32'b00000000000000000101001000111101; // input=-0.873046875, output=0.642494743009
			11'd1248: out = 32'b00000000000000000101000111011011; // input=-0.876953125, output=0.63949652811
			11'd1249: out = 32'b00000000000000000101000101111000; // input=-0.880859375, output=0.63648855528
			11'd1250: out = 32'b00000000000000000101000100010110; // input=-0.884765625, output=0.633470870418
			11'd1251: out = 32'b00000000000000000101000010110010; // input=-0.888671875, output=0.63044351957
			11'd1252: out = 32'b00000000000000000101000001001111; // input=-0.892578125, output=0.62740654893
			11'd1253: out = 32'b00000000000000000100111111101011; // input=-0.896484375, output=0.624360004837
			11'd1254: out = 32'b00000000000000000100111110000111; // input=-0.900390625, output=0.621303933779
			11'd1255: out = 32'b00000000000000000100111100100010; // input=-0.904296875, output=0.618238382388
			11'd1256: out = 32'b00000000000000000100111010111110; // input=-0.908203125, output=0.615163397439
			11'd1257: out = 32'b00000000000000000100111001011001; // input=-0.912109375, output=0.612079025854
			11'd1258: out = 32'b00000000000000000100110111110011; // input=-0.916015625, output=0.608985314696
			11'd1259: out = 32'b00000000000000000100110110001110; // input=-0.919921875, output=0.605882311171
			11'd1260: out = 32'b00000000000000000100110100101000; // input=-0.923828125, output=0.602770062628
			11'd1261: out = 32'b00000000000000000100110011000001; // input=-0.927734375, output=0.599648616555
			11'd1262: out = 32'b00000000000000000100110001011011; // input=-0.931640625, output=0.596518020582
			11'd1263: out = 32'b00000000000000000100101111110100; // input=-0.935546875, output=0.593378322478
			11'd1264: out = 32'b00000000000000000100101110001101; // input=-0.939453125, output=0.590229570151
			11'd1265: out = 32'b00000000000000000100101100100101; // input=-0.943359375, output=0.587071811646
			11'd1266: out = 32'b00000000000000000100101010111101; // input=-0.947265625, output=0.583905095149
			11'd1267: out = 32'b00000000000000000100101001010101; // input=-0.951171875, output=0.580729468977
			11'd1268: out = 32'b00000000000000000100100111101101; // input=-0.955078125, output=0.577544981589
			11'd1269: out = 32'b00000000000000000100100110000100; // input=-0.958984375, output=0.574351681575
			11'd1270: out = 32'b00000000000000000100100100011011; // input=-0.962890625, output=0.571149617661
			11'd1271: out = 32'b00000000000000000100100010110010; // input=-0.966796875, output=0.567938838706
			11'd1272: out = 32'b00000000000000000100100001001001; // input=-0.970703125, output=0.564719393703
			11'd1273: out = 32'b00000000000000000100011111011111; // input=-0.974609375, output=0.561491331777
			11'd1274: out = 32'b00000000000000000100011101110101; // input=-0.978515625, output=0.558254702185
			11'd1275: out = 32'b00000000000000000100011100001011; // input=-0.982421875, output=0.555009554312
			11'd1276: out = 32'b00000000000000000100011010100000; // input=-0.986328125, output=0.551755937677
			11'd1277: out = 32'b00000000000000000100011000110101; // input=-0.990234375, output=0.548493901924
			11'd1278: out = 32'b00000000000000000100010111001010; // input=-0.994140625, output=0.54522349683
			11'd1279: out = 32'b00000000000000000100010101011110; // input=-0.998046875, output=0.541944772296
			11'd1280: out = 32'b00000000000000000100010011110011; // input=-1.001953125, output=0.538657778351
			11'd1281: out = 32'b00000000000000000100010010000111; // input=-1.005859375, output=0.535362565152
			11'd1282: out = 32'b00000000000000000100010000011011; // input=-1.009765625, output=0.532059182978
			11'd1283: out = 32'b00000000000000000100001110101110; // input=-1.013671875, output=0.528747682236
			11'd1284: out = 32'b00000000000000000100001101000001; // input=-1.017578125, output=0.525428113455
			11'd1285: out = 32'b00000000000000000100001011010100; // input=-1.021484375, output=0.522100527287
			11'd1286: out = 32'b00000000000000000100001001100111; // input=-1.025390625, output=0.518764974507
			11'd1287: out = 32'b00000000000000000100000111111001; // input=-1.029296875, output=0.515421506013
			11'd1288: out = 32'b00000000000000000100000110001100; // input=-1.033203125, output=0.51207017282
			11'd1289: out = 32'b00000000000000000100000100011101; // input=-1.037109375, output=0.508711026066
			11'd1290: out = 32'b00000000000000000100000010101111; // input=-1.041015625, output=0.505344117008
			11'd1291: out = 32'b00000000000000000100000001000001; // input=-1.044921875, output=0.501969497021
			11'd1292: out = 32'b00000000000000000011111111010010; // input=-1.048828125, output=0.498587217597
			11'd1293: out = 32'b00000000000000000011111101100011; // input=-1.052734375, output=0.495197330345
			11'd1294: out = 32'b00000000000000000011111011110011; // input=-1.056640625, output=0.491799886991
			11'd1295: out = 32'b00000000000000000011111010000100; // input=-1.060546875, output=0.488394939376
			11'd1296: out = 32'b00000000000000000011111000010100; // input=-1.064453125, output=0.484982539455
			11'd1297: out = 32'b00000000000000000011110110100100; // input=-1.068359375, output=0.481562739297
			11'd1298: out = 32'b00000000000000000011110100110100; // input=-1.072265625, output=0.478135591084
			11'd1299: out = 32'b00000000000000000011110011000011; // input=-1.076171875, output=0.474701147111
			11'd1300: out = 32'b00000000000000000011110001010010; // input=-1.080078125, output=0.471259459782
			11'd1301: out = 32'b00000000000000000011101111100001; // input=-1.083984375, output=0.467810581613
			11'd1302: out = 32'b00000000000000000011101101110000; // input=-1.087890625, output=0.464354565231
			11'd1303: out = 32'b00000000000000000011101011111110; // input=-1.091796875, output=0.460891463369
			11'd1304: out = 32'b00000000000000000011101010001101; // input=-1.095703125, output=0.45742132887
			11'd1305: out = 32'b00000000000000000011101000011011; // input=-1.099609375, output=0.453944214685
			11'd1306: out = 32'b00000000000000000011100110101001; // input=-1.103515625, output=0.45046017387
			11'd1307: out = 32'b00000000000000000011100100110110; // input=-1.107421875, output=0.446969259586
			11'd1308: out = 32'b00000000000000000011100011000100; // input=-1.111328125, output=0.443471525102
			11'd1309: out = 32'b00000000000000000011100001010001; // input=-1.115234375, output=0.439967023787
			11'd1310: out = 32'b00000000000000000011011111011110; // input=-1.119140625, output=0.436455809118
			11'd1311: out = 32'b00000000000000000011011101101011; // input=-1.123046875, output=0.432937934669
			11'd1312: out = 32'b00000000000000000011011011110111; // input=-1.126953125, output=0.429413454121
			11'd1313: out = 32'b00000000000000000011011010000011; // input=-1.130859375, output=0.425882421251
			11'd1314: out = 32'b00000000000000000011011000001111; // input=-1.134765625, output=0.42234488994
			11'd1315: out = 32'b00000000000000000011010110011011; // input=-1.138671875, output=0.418800914165
			11'd1316: out = 32'b00000000000000000011010100100111; // input=-1.142578125, output=0.415250548003
			11'd1317: out = 32'b00000000000000000011010010110010; // input=-1.146484375, output=0.411693845629
			11'd1318: out = 32'b00000000000000000011010000111110; // input=-1.150390625, output=0.408130861314
			11'd1319: out = 32'b00000000000000000011001111001001; // input=-1.154296875, output=0.404561649424
			11'd1320: out = 32'b00000000000000000011001101010100; // input=-1.158203125, output=0.40098626442
			11'd1321: out = 32'b00000000000000000011001011011110; // input=-1.162109375, output=0.39740476086
			11'd1322: out = 32'b00000000000000000011001001101001; // input=-1.166015625, output=0.393817193392
			11'd1323: out = 32'b00000000000000000011000111110011; // input=-1.169921875, output=0.390223616758
			11'd1324: out = 32'b00000000000000000011000101111101; // input=-1.173828125, output=0.386624085792
			11'd1325: out = 32'b00000000000000000011000100000111; // input=-1.177734375, output=0.383018655418
			11'd1326: out = 32'b00000000000000000011000010010000; // input=-1.181640625, output=0.37940738065
			11'd1327: out = 32'b00000000000000000011000000011010; // input=-1.185546875, output=0.375790316593
			11'd1328: out = 32'b00000000000000000010111110100011; // input=-1.189453125, output=0.372167518438
			11'd1329: out = 32'b00000000000000000010111100101100; // input=-1.193359375, output=0.368539041464
			11'd1330: out = 32'b00000000000000000010111010110101; // input=-1.197265625, output=0.364904941038
			11'd1331: out = 32'b00000000000000000010111000111110; // input=-1.201171875, output=0.361265272612
			11'd1332: out = 32'b00000000000000000010110111000110; // input=-1.205078125, output=0.357620091721
			11'd1333: out = 32'b00000000000000000010110101001111; // input=-1.208984375, output=0.353969453989
			11'd1334: out = 32'b00000000000000000010110011010111; // input=-1.212890625, output=0.350313415118
			11'd1335: out = 32'b00000000000000000010110001011111; // input=-1.216796875, output=0.346652030895
			11'd1336: out = 32'b00000000000000000010101111100111; // input=-1.220703125, output=0.342985357189
			11'd1337: out = 32'b00000000000000000010101101101111; // input=-1.224609375, output=0.339313449948
			11'd1338: out = 32'b00000000000000000010101011110110; // input=-1.228515625, output=0.335636365202
			11'd1339: out = 32'b00000000000000000010101001111101; // input=-1.232421875, output=0.331954159057
			11'd1340: out = 32'b00000000000000000010101000000101; // input=-1.236328125, output=0.328266887701
			11'd1341: out = 32'b00000000000000000010100110001100; // input=-1.240234375, output=0.324574607395
			11'd1342: out = 32'b00000000000000000010100100010011; // input=-1.244140625, output=0.320877374481
			11'd1343: out = 32'b00000000000000000010100010011001; // input=-1.248046875, output=0.317175245372
			11'd1344: out = 32'b00000000000000000010100000100000; // input=-1.251953125, output=0.31346827656
			11'd1345: out = 32'b00000000000000000010011110100110; // input=-1.255859375, output=0.309756524607
			11'd1346: out = 32'b00000000000000000010011100101100; // input=-1.259765625, output=0.306040046151
			11'd1347: out = 32'b00000000000000000010011010110010; // input=-1.263671875, output=0.3023188979
			11'd1348: out = 32'b00000000000000000010011000111000; // input=-1.267578125, output=0.298593136635
			11'd1349: out = 32'b00000000000000000010010110111110; // input=-1.271484375, output=0.294862819205
			11'd1350: out = 32'b00000000000000000010010101000100; // input=-1.275390625, output=0.291128002532
			11'd1351: out = 32'b00000000000000000010010011001001; // input=-1.279296875, output=0.287388743604
			11'd1352: out = 32'b00000000000000000010010001001110; // input=-1.283203125, output=0.283645099478
			11'd1353: out = 32'b00000000000000000010001111010100; // input=-1.287109375, output=0.279897127276
			11'd1354: out = 32'b00000000000000000010001101011001; // input=-1.291015625, output=0.276144884188
			11'd1355: out = 32'b00000000000000000010001011011110; // input=-1.294921875, output=0.272388427469
			11'd1356: out = 32'b00000000000000000010001001100010; // input=-1.298828125, output=0.268627814438
			11'd1357: out = 32'b00000000000000000010000111100111; // input=-1.302734375, output=0.264863102477
			11'd1358: out = 32'b00000000000000000010000101101100; // input=-1.306640625, output=0.26109434903
			11'd1359: out = 32'b00000000000000000010000011110000; // input=-1.310546875, output=0.257321611606
			11'd1360: out = 32'b00000000000000000010000001110100; // input=-1.314453125, output=0.25354494777
			11'd1361: out = 32'b00000000000000000001111111111000; // input=-1.318359375, output=0.24976441515
			11'd1362: out = 32'b00000000000000000001111101111100; // input=-1.322265625, output=0.245980071432
			11'd1363: out = 32'b00000000000000000001111100000000; // input=-1.326171875, output=0.242191974361
			11'd1364: out = 32'b00000000000000000001111010000100; // input=-1.330078125, output=0.238400181739
			11'd1365: out = 32'b00000000000000000001111000001000; // input=-1.333984375, output=0.234604751423
			11'd1366: out = 32'b00000000000000000001110110001011; // input=-1.337890625, output=0.230805741327
			11'd1367: out = 32'b00000000000000000001110100001110; // input=-1.341796875, output=0.22700320942
			11'd1368: out = 32'b00000000000000000001110010010010; // input=-1.345703125, output=0.223197213723
			11'd1369: out = 32'b00000000000000000001110000010101; // input=-1.349609375, output=0.219387812311
			11'd1370: out = 32'b00000000000000000001101110011000; // input=-1.353515625, output=0.215575063311
			11'd1371: out = 32'b00000000000000000001101100011011; // input=-1.357421875, output=0.211759024901
			11'd1372: out = 32'b00000000000000000001101010011110; // input=-1.361328125, output=0.207939755308
			11'd1373: out = 32'b00000000000000000001101000100001; // input=-1.365234375, output=0.204117312811
			11'd1374: out = 32'b00000000000000000001100110100011; // input=-1.369140625, output=0.200291755735
			11'd1375: out = 32'b00000000000000000001100100100110; // input=-1.373046875, output=0.196463142453
			11'd1376: out = 32'b00000000000000000001100010101000; // input=-1.376953125, output=0.192631531385
			11'd1377: out = 32'b00000000000000000001100000101010; // input=-1.380859375, output=0.188796980997
			11'd1378: out = 32'b00000000000000000001011110101101; // input=-1.384765625, output=0.184959549799
			11'd1379: out = 32'b00000000000000000001011100101111; // input=-1.388671875, output=0.181119296346
			11'd1380: out = 32'b00000000000000000001011010110001; // input=-1.392578125, output=0.177276279236
			11'd1381: out = 32'b00000000000000000001011000110011; // input=-1.396484375, output=0.173430557107
			11'd1382: out = 32'b00000000000000000001010110110101; // input=-1.400390625, output=0.169582188642
			11'd1383: out = 32'b00000000000000000001010100110111; // input=-1.404296875, output=0.165731232561
			11'd1384: out = 32'b00000000000000000001010010111000; // input=-1.408203125, output=0.161877747625
			11'd1385: out = 32'b00000000000000000001010000111010; // input=-1.412109375, output=0.158021792634
			11'd1386: out = 32'b00000000000000000001001110111100; // input=-1.416015625, output=0.154163426425
			11'd1387: out = 32'b00000000000000000001001100111101; // input=-1.419921875, output=0.150302707872
			11'd1388: out = 32'b00000000000000000001001010111111; // input=-1.423828125, output=0.146439695884
			11'd1389: out = 32'b00000000000000000001001001000000; // input=-1.427734375, output=0.142574449407
			11'd1390: out = 32'b00000000000000000001000111000001; // input=-1.431640625, output=0.138707027419
			11'd1391: out = 32'b00000000000000000001000101000010; // input=-1.435546875, output=0.134837488933
			11'd1392: out = 32'b00000000000000000001000011000011; // input=-1.439453125, output=0.130965892992
			11'd1393: out = 32'b00000000000000000001000001000101; // input=-1.443359375, output=0.127092298673
			11'd1394: out = 32'b00000000000000000000111111000110; // input=-1.447265625, output=0.123216765082
			11'd1395: out = 32'b00000000000000000000111101000111; // input=-1.451171875, output=0.119339351355
			11'd1396: out = 32'b00000000000000000000111011000111; // input=-1.455078125, output=0.115460116656
			11'd1397: out = 32'b00000000000000000000111001001000; // input=-1.458984375, output=0.111579120177
			11'd1398: out = 32'b00000000000000000000110111001001; // input=-1.462890625, output=0.107696421139
			11'd1399: out = 32'b00000000000000000000110101001010; // input=-1.466796875, output=0.103812078785
			11'd1400: out = 32'b00000000000000000000110011001010; // input=-1.470703125, output=0.0999261523872
			11'd1401: out = 32'b00000000000000000000110001001011; // input=-1.474609375, output=0.0960387012391
			11'd1402: out = 32'b00000000000000000000101111001100; // input=-1.478515625, output=0.0921497846586
			11'd1403: out = 32'b00000000000000000000101101001100; // input=-1.482421875, output=0.0882594619857
			11'd1404: out = 32'b00000000000000000000101011001101; // input=-1.486328125, output=0.084367792582
			11'd1405: out = 32'b00000000000000000000101001001101; // input=-1.490234375, output=0.0804748358296
			11'd1406: out = 32'b00000000000000000000100111001101; // input=-1.494140625, output=0.0765806511302
			11'd1407: out = 32'b00000000000000000000100101001110; // input=-1.498046875, output=0.0726852979043
			11'd1408: out = 32'b00000000000000000000100011001110; // input=-1.501953125, output=0.0687888355902
			11'd1409: out = 32'b00000000000000000000100001001110; // input=-1.505859375, output=0.0648913236431
			11'd1410: out = 32'b00000000000000000000011111001111; // input=-1.509765625, output=0.0609928215342
			11'd1411: out = 32'b00000000000000000000011101001111; // input=-1.513671875, output=0.0570933887499
			11'd1412: out = 32'b00000000000000000000011011001111; // input=-1.517578125, output=0.0531930847907
			11'd1413: out = 32'b00000000000000000000011001001111; // input=-1.521484375, output=0.0492919691706
			11'd1414: out = 32'b00000000000000000000010111001111; // input=-1.525390625, output=0.0453901014156
			11'd1415: out = 32'b00000000000000000000010101001111; // input=-1.529296875, output=0.0414875410635
			11'd1416: out = 32'b00000000000000000000010011010000; // input=-1.533203125, output=0.0375843476626
			11'd1417: out = 32'b00000000000000000000010001010000; // input=-1.537109375, output=0.0336805807707
			11'd1418: out = 32'b00000000000000000000001111010000; // input=-1.541015625, output=0.0297762999547
			11'd1419: out = 32'b00000000000000000000001101010000; // input=-1.544921875, output=0.0258715647889
			11'd1420: out = 32'b00000000000000000000001011010000; // input=-1.548828125, output=0.0219664348549
			11'd1421: out = 32'b00000000000000000000001001010000; // input=-1.552734375, output=0.0180609697401
			11'd1422: out = 32'b00000000000000000000000111010000; // input=-1.556640625, output=0.0141552290372
			11'd1423: out = 32'b00000000000000000000000101010000; // input=-1.560546875, output=0.0102492723429
			11'd1424: out = 32'b00000000000000000000000011010000; // input=-1.564453125, output=0.00634315925725
			11'd1425: out = 32'b00000000000000000000000001010000; // input=-1.568359375, output=0.00243694938283
			11'd1426: out = 32'b10000000000000000000000000110000; // input=-1.572265625, output=-0.00146929767644
			11'd1427: out = 32'b10000000000000000000000010110000; // input=-1.576171875, output=-0.00537552231604
			11'd1428: out = 32'b10000000000000000000000100110000; // input=-1.580078125, output=-0.00928166493177
			11'd1429: out = 32'b10000000000000000000000110110000; // input=-1.583984375, output=-0.0131876659207
			11'd1430: out = 32'b10000000000000000000001000110000; // input=-1.587890625, output=-0.0170934656821
			11'd1431: out = 32'b10000000000000000000001010110000; // input=-1.591796875, output=-0.0209990046183
			11'd1432: out = 32'b10000000000000000000001100110000; // input=-1.595703125, output=-0.0249042231354
			11'd1433: out = 32'b10000000000000000000001110110000; // input=-1.599609375, output=-0.0288090616448
			11'd1434: out = 32'b10000000000000000000010000110000; // input=-1.603515625, output=-0.0327134605633
			11'd1435: out = 32'b10000000000000000000010010110000; // input=-1.607421875, output=-0.0366173603147
			11'd1436: out = 32'b10000000000000000000010100110000; // input=-1.611328125, output=-0.0405207013302
			11'd1437: out = 32'b10000000000000000000010110110000; // input=-1.615234375, output=-0.0444234240496
			11'd1438: out = 32'b10000000000000000000011000110000; // input=-1.619140625, output=-0.0483254689223
			11'd1439: out = 32'b10000000000000000000011010101111; // input=-1.623046875, output=-0.0522267764077
			11'd1440: out = 32'b10000000000000000000011100101111; // input=-1.626953125, output=-0.0561272869768
			11'd1441: out = 32'b10000000000000000000011110101111; // input=-1.630859375, output=-0.0600269411126
			11'd1442: out = 32'b10000000000000000000100000101111; // input=-1.634765625, output=-0.0639256793111
			11'd1443: out = 32'b10000000000000000000100010101110; // input=-1.638671875, output=-0.0678234420824
			11'd1444: out = 32'b10000000000000000000100100101110; // input=-1.642578125, output=-0.0717201699514
			11'd1445: out = 32'b10000000000000000000100110101110; // input=-1.646484375, output=-0.0756158034588
			11'd1446: out = 32'b10000000000000000000101000101101; // input=-1.650390625, output=-0.0795102831621
			11'd1447: out = 32'b10000000000000000000101010101101; // input=-1.654296875, output=-0.0834035496363
			11'd1448: out = 32'b10000000000000000000101100101101; // input=-1.658203125, output=-0.087295543475
			11'd1449: out = 32'b10000000000000000000101110101100; // input=-1.662109375, output=-0.0911862052911
			11'd1450: out = 32'b10000000000000000000110000101011; // input=-1.666015625, output=-0.0950754757179
			11'd1451: out = 32'b10000000000000000000110010101011; // input=-1.669921875, output=-0.0989632954099
			11'd1452: out = 32'b10000000000000000000110100101010; // input=-1.673828125, output=-0.102849605044
			11'd1453: out = 32'b10000000000000000000110110101001; // input=-1.677734375, output=-0.106734345319
			11'd1454: out = 32'b10000000000000000000111000101001; // input=-1.681640625, output=-0.11061745696
			11'd1455: out = 32'b10000000000000000000111010101000; // input=-1.685546875, output=-0.114498880714
			11'd1456: out = 32'b10000000000000000000111100100111; // input=-1.689453125, output=-0.118378557356
			11'd1457: out = 32'b10000000000000000000111110100110; // input=-1.693359375, output=-0.122256427688
			11'd1458: out = 32'b10000000000000000001000000100101; // input=-1.697265625, output=-0.126132432536
			11'd1459: out = 32'b10000000000000000001000010100100; // input=-1.701171875, output=-0.130006512759
			11'd1460: out = 32'b10000000000000000001000100100011; // input=-1.705078125, output=-0.133878609242
			11'd1461: out = 32'b10000000000000000001000110100010; // input=-1.708984375, output=-0.137748662903
			11'd1462: out = 32'b10000000000000000001001000100000; // input=-1.712890625, output=-0.141616614688
			11'd1463: out = 32'b10000000000000000001001010011111; // input=-1.716796875, output=-0.145482405578
			11'd1464: out = 32'b10000000000000000001001100011110; // input=-1.720703125, output=-0.149345976585
			11'd1465: out = 32'b10000000000000000001001110011100; // input=-1.724609375, output=-0.153207268757
			11'd1466: out = 32'b10000000000000000001010000011011; // input=-1.728515625, output=-0.157066223174
			11'd1467: out = 32'b10000000000000000001010010011001; // input=-1.732421875, output=-0.160922780954
			11'd1468: out = 32'b10000000000000000001010100010111; // input=-1.736328125, output=-0.164776883251
			11'd1469: out = 32'b10000000000000000001010110010110; // input=-1.740234375, output=-0.168628471254
			11'd1470: out = 32'b10000000000000000001011000010100; // input=-1.744140625, output=-0.172477486195
			11'd1471: out = 32'b10000000000000000001011010010010; // input=-1.748046875, output=-0.176323869342
			11'd1472: out = 32'b10000000000000000001011100010000; // input=-1.751953125, output=-0.180167562003
			11'd1473: out = 32'b10000000000000000001011110001110; // input=-1.755859375, output=-0.184008505529
			11'd1474: out = 32'b10000000000000000001100000001011; // input=-1.759765625, output=-0.187846641311
			11'd1475: out = 32'b10000000000000000001100010001001; // input=-1.763671875, output=-0.191681910785
			11'd1476: out = 32'b10000000000000000001100100000111; // input=-1.767578125, output=-0.195514255429
			11'd1477: out = 32'b10000000000000000001100110000100; // input=-1.771484375, output=-0.199343616766
			11'd1478: out = 32'b10000000000000000001101000000001; // input=-1.775390625, output=-0.203169936364
			11'd1479: out = 32'b10000000000000000001101001111111; // input=-1.779296875, output=-0.206993155839
			11'd1480: out = 32'b10000000000000000001101011111100; // input=-1.783203125, output=-0.210813216853
			11'd1481: out = 32'b10000000000000000001101101111001; // input=-1.787109375, output=-0.214630061117
			11'd1482: out = 32'b10000000000000000001101111110110; // input=-1.791015625, output=-0.218443630391
			11'd1483: out = 32'b10000000000000000001110001110011; // input=-1.794921875, output=-0.222253866483
			11'd1484: out = 32'b10000000000000000001110011110000; // input=-1.798828125, output=-0.226060711255
			11'd1485: out = 32'b10000000000000000001110101101100; // input=-1.802734375, output=-0.229864106618
			11'd1486: out = 32'b10000000000000000001110111101001; // input=-1.806640625, output=-0.233663994538
			11'd1487: out = 32'b10000000000000000001111001100101; // input=-1.810546875, output=-0.237460317033
			11'd1488: out = 32'b10000000000000000001111011100001; // input=-1.814453125, output=-0.241253016175
			11'd1489: out = 32'b10000000000000000001111101011110; // input=-1.818359375, output=-0.245042034094
			11'd1490: out = 32'b10000000000000000001111111011010; // input=-1.822265625, output=-0.248827312972
			11'd1491: out = 32'b10000000000000000010000001010101; // input=-1.826171875, output=-0.252608795052
			11'd1492: out = 32'b10000000000000000010000011010001; // input=-1.830078125, output=-0.256386422632
			11'd1493: out = 32'b10000000000000000010000101001101; // input=-1.833984375, output=-0.260160138071
			11'd1494: out = 32'b10000000000000000010000111001000; // input=-1.837890625, output=-0.263929883786
			11'd1495: out = 32'b10000000000000000010001001000100; // input=-1.841796875, output=-0.267695602256
			11'd1496: out = 32'b10000000000000000010001010111111; // input=-1.845703125, output=-0.271457236021
			11'd1497: out = 32'b10000000000000000010001100111010; // input=-1.849609375, output=-0.275214727682
			11'd1498: out = 32'b10000000000000000010001110110101; // input=-1.853515625, output=-0.278968019905
			11'd1499: out = 32'b10000000000000000010010000110000; // input=-1.857421875, output=-0.282717055419
			11'd1500: out = 32'b10000000000000000010010010101011; // input=-1.861328125, output=-0.286461777019
			11'd1501: out = 32'b10000000000000000010010100100101; // input=-1.865234375, output=-0.290202127564
			11'd1502: out = 32'b10000000000000000010010110100000; // input=-1.869140625, output=-0.293938049982
			11'd1503: out = 32'b10000000000000000010011000011010; // input=-1.873046875, output=-0.297669487267
			11'd1504: out = 32'b10000000000000000010011010010100; // input=-1.876953125, output=-0.301396382482
			11'd1505: out = 32'b10000000000000000010011100001110; // input=-1.880859375, output=-0.305118678759
			11'd1506: out = 32'b10000000000000000010011110001000; // input=-1.884765625, output=-0.308836319301
			11'd1507: out = 32'b10000000000000000010100000000010; // input=-1.888671875, output=-0.31254924738
			11'd1508: out = 32'b10000000000000000010100001111011; // input=-1.892578125, output=-0.316257406342
			11'd1509: out = 32'b10000000000000000010100011110100; // input=-1.896484375, output=-0.319960739605
			11'd1510: out = 32'b10000000000000000010100101101110; // input=-1.900390625, output=-0.323659190661
			11'd1511: out = 32'b10000000000000000010100111100111; // input=-1.904296875, output=-0.327352703076
			11'd1512: out = 32'b10000000000000000010101001100000; // input=-1.908203125, output=-0.331041220491
			11'd1513: out = 32'b10000000000000000010101011011000; // input=-1.912109375, output=-0.334724686625
			11'd1514: out = 32'b10000000000000000010101101010001; // input=-1.916015625, output=-0.338403045272
			11'd1515: out = 32'b10000000000000000010101111001001; // input=-1.919921875, output=-0.342076240304
			11'd1516: out = 32'b10000000000000000010110001000001; // input=-1.923828125, output=-0.345744215674
			11'd1517: out = 32'b10000000000000000010110010111001; // input=-1.927734375, output=-0.349406915413
			11'd1518: out = 32'b10000000000000000010110100110001; // input=-1.931640625, output=-0.353064283632
			11'd1519: out = 32'b10000000000000000010110110101001; // input=-1.935546875, output=-0.356716264525
			11'd1520: out = 32'b10000000000000000010111000100000; // input=-1.939453125, output=-0.360362802366
			11'd1521: out = 32'b10000000000000000010111010011000; // input=-1.943359375, output=-0.364003841514
			11'd1522: out = 32'b10000000000000000010111100001111; // input=-1.947265625, output=-0.367639326412
			11'd1523: out = 32'b10000000000000000010111110000110; // input=-1.951171875, output=-0.371269201585
			11'd1524: out = 32'b10000000000000000010111111111101; // input=-1.955078125, output=-0.374893411648
			11'd1525: out = 32'b10000000000000000011000001110011; // input=-1.958984375, output=-0.378511901298
			11'd1526: out = 32'b10000000000000000011000011101001; // input=-1.962890625, output=-0.382124615322
			11'd1527: out = 32'b10000000000000000011000101100000; // input=-1.966796875, output=-0.385731498595
			11'd1528: out = 32'b10000000000000000011000111010110; // input=-1.970703125, output=-0.38933249608
			11'd1529: out = 32'b10000000000000000011001001001011; // input=-1.974609375, output=-0.392927552829
			11'd1530: out = 32'b10000000000000000011001011000001; // input=-1.978515625, output=-0.396516613988
			11'd1531: out = 32'b10000000000000000011001100110110; // input=-1.982421875, output=-0.400099624791
			11'd1532: out = 32'b10000000000000000011001110101100; // input=-1.986328125, output=-0.403676530566
			11'd1533: out = 32'b10000000000000000011010000100001; // input=-1.990234375, output=-0.407247276734
			11'd1534: out = 32'b10000000000000000011010010010101; // input=-1.994140625, output=-0.41081180881
			11'd1535: out = 32'b10000000000000000011010100001010; // input=-1.998046875, output=-0.414370072403
			11'd1536: out = 32'b10000000000000000011010101111110; // input=-2.001953125, output=-0.417922013218
			11'd1537: out = 32'b10000000000000000011010111110011; // input=-2.005859375, output=-0.421467577057
			11'd1538: out = 32'b10000000000000000011011001100111; // input=-2.009765625, output=-0.42500670982
			11'd1539: out = 32'b10000000000000000011011011011010; // input=-2.013671875, output=-0.428539357504
			11'd1540: out = 32'b10000000000000000011011101001110; // input=-2.017578125, output=-0.432065466204
			11'd1541: out = 32'b10000000000000000011011111000001; // input=-2.021484375, output=-0.435584982116
			11'd1542: out = 32'b10000000000000000011100000110100; // input=-2.025390625, output=-0.439097851538
			11'd1543: out = 32'b10000000000000000011100010100111; // input=-2.029296875, output=-0.442604020867
			11'd1544: out = 32'b10000000000000000011100100011010; // input=-2.033203125, output=-0.446103436603
			11'd1545: out = 32'b10000000000000000011100110001100; // input=-2.037109375, output=-0.449596045349
			11'd1546: out = 32'b10000000000000000011100111111111; // input=-2.041015625, output=-0.453081793813
			11'd1547: out = 32'b10000000000000000011101001110001; // input=-2.044921875, output=-0.456560628806
			11'd1548: out = 32'b10000000000000000011101011100010; // input=-2.048828125, output=-0.460032497246
			11'd1549: out = 32'b10000000000000000011101101010100; // input=-2.052734375, output=-0.463497346155
			11'd1550: out = 32'b10000000000000000011101111000101; // input=-2.056640625, output=-0.466955122666
			11'd1551: out = 32'b10000000000000000011110000110110; // input=-2.060546875, output=-0.470405774016
			11'd1552: out = 32'b10000000000000000011110010100111; // input=-2.064453125, output=-0.473849247552
			11'd1553: out = 32'b10000000000000000011110100011000; // input=-2.068359375, output=-0.477285490732
			11'd1554: out = 32'b10000000000000000011110110001000; // input=-2.072265625, output=-0.480714451123
			11'd1555: out = 32'b10000000000000000011110111111000; // input=-2.076171875, output=-0.484136076402
			11'd1556: out = 32'b10000000000000000011111001101000; // input=-2.080078125, output=-0.487550314361
			11'd1557: out = 32'b10000000000000000011111011011000; // input=-2.083984375, output=-0.490957112901
			11'd1558: out = 32'b10000000000000000011111101000111; // input=-2.087890625, output=-0.49435642004
			11'd1559: out = 32'b10000000000000000011111110110110; // input=-2.091796875, output=-0.497748183909
			11'd1560: out = 32'b10000000000000000100000000100101; // input=-2.095703125, output=-0.501132352752
			11'd1561: out = 32'b10000000000000000100000010010100; // input=-2.099609375, output=-0.504508874933
			11'd1562: out = 32'b10000000000000000100000100000010; // input=-2.103515625, output=-0.507877698929
			11'd1563: out = 32'b10000000000000000100000101110000; // input=-2.107421875, output=-0.511238773335
			11'd1564: out = 32'b10000000000000000100000111011110; // input=-2.111328125, output=-0.514592046868
			11'd1565: out = 32'b10000000000000000100001001001100; // input=-2.115234375, output=-0.517937468358
			11'd1566: out = 32'b10000000000000000100001010111001; // input=-2.119140625, output=-0.52127498676
			11'd1567: out = 32'b10000000000000000100001100100110; // input=-2.123046875, output=-0.524604551148
			11'd1568: out = 32'b10000000000000000100001110010011; // input=-2.126953125, output=-0.527926110715
			11'd1569: out = 32'b10000000000000000100010000000000; // input=-2.130859375, output=-0.531239614779
			11'd1570: out = 32'b10000000000000000100010001101100; // input=-2.134765625, output=-0.53454501278
			11'd1571: out = 32'b10000000000000000100010011011000; // input=-2.138671875, output=-0.537842254283
			11'd1572: out = 32'b10000000000000000100010101000100; // input=-2.142578125, output=-0.541131288974
			11'd1573: out = 32'b10000000000000000100010110101111; // input=-2.146484375, output=-0.544412066667
			11'd1574: out = 32'b10000000000000000100011000011011; // input=-2.150390625, output=-0.547684537302
			11'd1575: out = 32'b10000000000000000100011010000101; // input=-2.154296875, output=-0.550948650945
			11'd1576: out = 32'b10000000000000000100011011110000; // input=-2.158203125, output=-0.554204357789
			11'd1577: out = 32'b10000000000000000100011101011011; // input=-2.162109375, output=-0.557451608157
			11'd1578: out = 32'b10000000000000000100011111000101; // input=-2.166015625, output=-0.560690352499
			11'd1579: out = 32'b10000000000000000100100000101111; // input=-2.169921875, output=-0.563920541396
			11'd1580: out = 32'b10000000000000000100100010011000; // input=-2.173828125, output=-0.567142125559
			11'd1581: out = 32'b10000000000000000100100100000001; // input=-2.177734375, output=-0.570355055831
			11'd1582: out = 32'b10000000000000000100100101101010; // input=-2.181640625, output=-0.573559283187
			11'd1583: out = 32'b10000000000000000100100111010011; // input=-2.185546875, output=-0.576754758734
			11'd1584: out = 32'b10000000000000000100101000111100; // input=-2.189453125, output=-0.579941433713
			11'd1585: out = 32'b10000000000000000100101010100100; // input=-2.193359375, output=-0.583119259499
			11'd1586: out = 32'b10000000000000000100101100001011; // input=-2.197265625, output=-0.586288187603
			11'd1587: out = 32'b10000000000000000100101101110011; // input=-2.201171875, output=-0.58944816967
			11'd1588: out = 32'b10000000000000000100101111011010; // input=-2.205078125, output=-0.592599157484
			11'd1589: out = 32'b10000000000000000100110001000001; // input=-2.208984375, output=-0.595741102963
			11'd1590: out = 32'b10000000000000000100110010101000; // input=-2.212890625, output=-0.598873958166
			11'd1591: out = 32'b10000000000000000100110100001110; // input=-2.216796875, output=-0.601997675289
			11'd1592: out = 32'b10000000000000000100110101110100; // input=-2.220703125, output=-0.605112206669
			11'd1593: out = 32'b10000000000000000100110111011010; // input=-2.224609375, output=-0.60821750478
			11'd1594: out = 32'b10000000000000000100111001000000; // input=-2.228515625, output=-0.611313522241
			11'd1595: out = 32'b10000000000000000100111010100101; // input=-2.232421875, output=-0.61440021181
			11'd1596: out = 32'b10000000000000000100111100001010; // input=-2.236328125, output=-0.617477526387
			11'd1597: out = 32'b10000000000000000100111101101110; // input=-2.240234375, output=-0.620545419017
			11'd1598: out = 32'b10000000000000000100111111010010; // input=-2.244140625, output=-0.623603842888
			11'd1599: out = 32'b10000000000000000101000000110110; // input=-2.248046875, output=-0.626652751331
			11'd1600: out = 32'b10000000000000000101000010011010; // input=-2.251953125, output=-0.629692097824
			11'd1601: out = 32'b10000000000000000101000011111101; // input=-2.255859375, output=-0.63272183599
			11'd1602: out = 32'b10000000000000000101000101100000; // input=-2.259765625, output=-0.635741919599
			11'd1603: out = 32'b10000000000000000101000111000011; // input=-2.263671875, output=-0.638752302569
			11'd1604: out = 32'b10000000000000000101001000100101; // input=-2.267578125, output=-0.641752938965
			11'd1605: out = 32'b10000000000000000101001010000111; // input=-2.271484375, output=-0.644743783001
			11'd1606: out = 32'b10000000000000000101001011101001; // input=-2.275390625, output=-0.647724789039
			11'd1607: out = 32'b10000000000000000101001101001010; // input=-2.279296875, output=-0.650695911595
			11'd1608: out = 32'b10000000000000000101001110101011; // input=-2.283203125, output=-0.653657105331
			11'd1609: out = 32'b10000000000000000101010000001100; // input=-2.287109375, output=-0.656608325064
			11'd1610: out = 32'b10000000000000000101010001101100; // input=-2.291015625, output=-0.659549525762
			11'd1611: out = 32'b10000000000000000101010011001100; // input=-2.294921875, output=-0.662480662545
			11'd1612: out = 32'b10000000000000000101010100101100; // input=-2.298828125, output=-0.665401690689
			11'd1613: out = 32'b10000000000000000101010110001011; // input=-2.302734375, output=-0.668312565622
			11'd1614: out = 32'b10000000000000000101010111101010; // input=-2.306640625, output=-0.671213242927
			11'd1615: out = 32'b10000000000000000101011001001001; // input=-2.310546875, output=-0.674103678343
			11'd1616: out = 32'b10000000000000000101011010100111; // input=-2.314453125, output=-0.676983827767
			11'd1617: out = 32'b10000000000000000101011100000101; // input=-2.318359375, output=-0.679853647251
			11'd1618: out = 32'b10000000000000000101011101100011; // input=-2.322265625, output=-0.682713093005
			11'd1619: out = 32'b10000000000000000101011111000000; // input=-2.326171875, output=-0.685562121397
			11'd1620: out = 32'b10000000000000000101100000011110; // input=-2.330078125, output=-0.688400688954
			11'd1621: out = 32'b10000000000000000101100001111010; // input=-2.333984375, output=-0.691228752363
			11'd1622: out = 32'b10000000000000000101100011010111; // input=-2.337890625, output=-0.694046268473
			11'd1623: out = 32'b10000000000000000101100100110010; // input=-2.341796875, output=-0.69685319429
			11'd1624: out = 32'b10000000000000000101100110001110; // input=-2.345703125, output=-0.699649486985
			11'd1625: out = 32'b10000000000000000101100111101001; // input=-2.349609375, output=-0.702435103889
			11'd1626: out = 32'b10000000000000000101101001000100; // input=-2.353515625, output=-0.705210002498
			11'd1627: out = 32'b10000000000000000101101010011111; // input=-2.357421875, output=-0.707974140471
			11'd1628: out = 32'b10000000000000000101101011111001; // input=-2.361328125, output=-0.710727475628
			11'd1629: out = 32'b10000000000000000101101101010011; // input=-2.365234375, output=-0.713469965959
			11'd1630: out = 32'b10000000000000000101101110101100; // input=-2.369140625, output=-0.716201569616
			11'd1631: out = 32'b10000000000000000101110000000110; // input=-2.373046875, output=-0.718922244918
			11'd1632: out = 32'b10000000000000000101110001011110; // input=-2.376953125, output=-0.721631950352
			11'd1633: out = 32'b10000000000000000101110010110111; // input=-2.380859375, output=-0.724330644569
			11'd1634: out = 32'b10000000000000000101110100001111; // input=-2.384765625, output=-0.727018286392
			11'd1635: out = 32'b10000000000000000101110101100111; // input=-2.388671875, output=-0.729694834811
			11'd1636: out = 32'b10000000000000000101110110111110; // input=-2.392578125, output=-0.732360248984
			11'd1637: out = 32'b10000000000000000101111000010101; // input=-2.396484375, output=-0.735014488241
			11'd1638: out = 32'b10000000000000000101111001101100; // input=-2.400390625, output=-0.737657512081
			11'd1639: out = 32'b10000000000000000101111011000010; // input=-2.404296875, output=-0.740289280175
			11'd1640: out = 32'b10000000000000000101111100011000; // input=-2.408203125, output=-0.742909752365
			11'd1641: out = 32'b10000000000000000101111101101101; // input=-2.412109375, output=-0.745518888667
			11'd1642: out = 32'b10000000000000000101111111000010; // input=-2.416015625, output=-0.748116649267
			11'd1643: out = 32'b10000000000000000110000000010111; // input=-2.419921875, output=-0.750702994528
			11'd1644: out = 32'b10000000000000000110000001101011; // input=-2.423828125, output=-0.753277884985
			11'd1645: out = 32'b10000000000000000110000010111111; // input=-2.427734375, output=-0.755841281348
			11'd1646: out = 32'b10000000000000000110000100010011; // input=-2.431640625, output=-0.758393144503
			11'd1647: out = 32'b10000000000000000110000101100110; // input=-2.435546875, output=-0.760933435512
			11'd1648: out = 32'b10000000000000000110000110111001; // input=-2.439453125, output=-0.763462115613
			11'd1649: out = 32'b10000000000000000110001000001100; // input=-2.443359375, output=-0.765979146221
			11'd1650: out = 32'b10000000000000000110001001011110; // input=-2.447265625, output=-0.76848448893
			11'd1651: out = 32'b10000000000000000110001010101111; // input=-2.451171875, output=-0.770978105511
			11'd1652: out = 32'b10000000000000000110001100000001; // input=-2.455078125, output=-0.773459957915
			11'd1653: out = 32'b10000000000000000110001101010010; // input=-2.458984375, output=-0.775930008271
			11'd1654: out = 32'b10000000000000000110001110100010; // input=-2.462890625, output=-0.77838821889
			11'd1655: out = 32'b10000000000000000110001111110010; // input=-2.466796875, output=-0.780834552263
			11'd1656: out = 32'b10000000000000000110010001000010; // input=-2.470703125, output=-0.783268971061
			11'd1657: out = 32'b10000000000000000110010010010010; // input=-2.474609375, output=-0.785691438138
			11'd1658: out = 32'b10000000000000000110010011100001; // input=-2.478515625, output=-0.78810191653
			11'd1659: out = 32'b10000000000000000110010100101111; // input=-2.482421875, output=-0.790500369457
			11'd1660: out = 32'b10000000000000000110010101111101; // input=-2.486328125, output=-0.792886760321
			11'd1661: out = 32'b10000000000000000110010111001011; // input=-2.490234375, output=-0.795261052708
			11'd1662: out = 32'b10000000000000000110011000011001; // input=-2.494140625, output=-0.797623210391
			11'd1663: out = 32'b10000000000000000110011001100110; // input=-2.498046875, output=-0.799973197324
			11'd1664: out = 32'b10000000000000000110011010110010; // input=-2.501953125, output=-0.802310977651
			11'd1665: out = 32'b10000000000000000110011011111110; // input=-2.505859375, output=-0.804636515699
			11'd1666: out = 32'b10000000000000000110011101001010; // input=-2.509765625, output=-0.806949775984
			11'd1667: out = 32'b10000000000000000110011110010110; // input=-2.513671875, output=-0.809250723208
			11'd1668: out = 32'b10000000000000000110011111100001; // input=-2.517578125, output=-0.811539322262
			11'd1669: out = 32'b10000000000000000110100000101011; // input=-2.521484375, output=-0.813815538224
			11'd1670: out = 32'b10000000000000000110100001110101; // input=-2.525390625, output=-0.816079336362
			11'd1671: out = 32'b10000000000000000110100010111111; // input=-2.529296875, output=-0.818330682134
			11'd1672: out = 32'b10000000000000000110100100001000; // input=-2.533203125, output=-0.820569541186
			11'd1673: out = 32'b10000000000000000110100101010001; // input=-2.537109375, output=-0.822795879357
			11'd1674: out = 32'b10000000000000000110100110011010; // input=-2.541015625, output=-0.825009662675
			11'd1675: out = 32'b10000000000000000110100111100010; // input=-2.544921875, output=-0.82721085736
			11'd1676: out = 32'b10000000000000000110101000101010; // input=-2.548828125, output=-0.829399429826
			11'd1677: out = 32'b10000000000000000110101001110001; // input=-2.552734375, output=-0.831575346677
			11'd1678: out = 32'b10000000000000000110101010111000; // input=-2.556640625, output=-0.833738574711
			11'd1679: out = 32'b10000000000000000110101011111110; // input=-2.560546875, output=-0.83588908092
			11'd1680: out = 32'b10000000000000000110101101000100; // input=-2.564453125, output=-0.83802683249
			11'd1681: out = 32'b10000000000000000110101110001010; // input=-2.568359375, output=-0.840151796802
			11'd1682: out = 32'b10000000000000000110101111001111; // input=-2.572265625, output=-0.842263941431
			11'd1683: out = 32'b10000000000000000110110000010100; // input=-2.576171875, output=-0.844363234149
			11'd1684: out = 32'b10000000000000000110110001011000; // input=-2.580078125, output=-0.846449642922
			11'd1685: out = 32'b10000000000000000110110010011100; // input=-2.583984375, output=-0.848523135916
			11'd1686: out = 32'b10000000000000000110110011100000; // input=-2.587890625, output=-0.85058368149
			11'd1687: out = 32'b10000000000000000110110100100011; // input=-2.591796875, output=-0.852631248204
			11'd1688: out = 32'b10000000000000000110110101100110; // input=-2.595703125, output=-0.854665804814
			11'd1689: out = 32'b10000000000000000110110110101000; // input=-2.599609375, output=-0.856687320275
			11'd1690: out = 32'b10000000000000000110110111101010; // input=-2.603515625, output=-0.858695763742
			11'd1691: out = 32'b10000000000000000110111000101011; // input=-2.607421875, output=-0.860691104568
			11'd1692: out = 32'b10000000000000000110111001101100; // input=-2.611328125, output=-0.862673312307
			11'd1693: out = 32'b10000000000000000110111010101101; // input=-2.615234375, output=-0.864642356712
			11'd1694: out = 32'b10000000000000000110111011101101; // input=-2.619140625, output=-0.866598207739
			11'd1695: out = 32'b10000000000000000110111100101100; // input=-2.623046875, output=-0.868540835543
			11'd1696: out = 32'b10000000000000000110111101101100; // input=-2.626953125, output=-0.870470210483
			11'd1697: out = 32'b10000000000000000110111110101010; // input=-2.630859375, output=-0.872386303118
			11'd1698: out = 32'b10000000000000000110111111101001; // input=-2.634765625, output=-0.874289084212
			11'd1699: out = 32'b10000000000000000111000000100111; // input=-2.638671875, output=-0.87617852473
			11'd1700: out = 32'b10000000000000000111000001100100; // input=-2.642578125, output=-0.878054595842
			11'd1701: out = 32'b10000000000000000111000010100001; // input=-2.646484375, output=-0.879917268921
			11'd1702: out = 32'b10000000000000000111000011011110; // input=-2.650390625, output=-0.881766515544
			11'd1703: out = 32'b10000000000000000111000100011010; // input=-2.654296875, output=-0.883602307496
			11'd1704: out = 32'b10000000000000000111000101010110; // input=-2.658203125, output=-0.885424616764
			11'd1705: out = 32'b10000000000000000111000110010001; // input=-2.662109375, output=-0.887233415541
			11'd1706: out = 32'b10000000000000000111000111001100; // input=-2.666015625, output=-0.889028676228
			11'd1707: out = 32'b10000000000000000111001000000110; // input=-2.669921875, output=-0.890810371432
			11'd1708: out = 32'b10000000000000000111001001000000; // input=-2.673828125, output=-0.892578473965
			11'd1709: out = 32'b10000000000000000111001001111010; // input=-2.677734375, output=-0.894332956848
			11'd1710: out = 32'b10000000000000000111001010110011; // input=-2.681640625, output=-0.896073793311
			11'd1711: out = 32'b10000000000000000111001011101011; // input=-2.685546875, output=-0.897800956791
			11'd1712: out = 32'b10000000000000000111001100100011; // input=-2.689453125, output=-0.899514420932
			11'd1713: out = 32'b10000000000000000111001101011011; // input=-2.693359375, output=-0.90121415959
			11'd1714: out = 32'b10000000000000000111001110010010; // input=-2.697265625, output=-0.902900146829
			11'd1715: out = 32'b10000000000000000111001111001001; // input=-2.701171875, output=-0.904572356923
			11'd1716: out = 32'b10000000000000000111001111111111; // input=-2.705078125, output=-0.906230764355
			11'd1717: out = 32'b10000000000000000111010000110101; // input=-2.708984375, output=-0.907875343821
			11'd1718: out = 32'b10000000000000000111010001101011; // input=-2.712890625, output=-0.909506070226
			11'd1719: out = 32'b10000000000000000111010010100000; // input=-2.716796875, output=-0.911122918687
			11'd1720: out = 32'b10000000000000000111010011010100; // input=-2.720703125, output=-0.912725864533
			11'd1721: out = 32'b10000000000000000111010100001000; // input=-2.724609375, output=-0.914314883306
			11'd1722: out = 32'b10000000000000000111010100111100; // input=-2.728515625, output=-0.915889950759
			11'd1723: out = 32'b10000000000000000111010101101111; // input=-2.732421875, output=-0.917451042858
			11'd1724: out = 32'b10000000000000000111010110100010; // input=-2.736328125, output=-0.918998135783
			11'd1725: out = 32'b10000000000000000111010111010100; // input=-2.740234375, output=-0.920531205927
			11'd1726: out = 32'b10000000000000000111011000000110; // input=-2.744140625, output=-0.922050229897
			11'd1727: out = 32'b10000000000000000111011000110111; // input=-2.748046875, output=-0.923555184515
			11'd1728: out = 32'b10000000000000000111011001101000; // input=-2.751953125, output=-0.925046046817
			11'd1729: out = 32'b10000000000000000111011010011000; // input=-2.755859375, output=-0.926522794055
			11'd1730: out = 32'b10000000000000000111011011001000; // input=-2.759765625, output=-0.927985403695
			11'd1731: out = 32'b10000000000000000111011011111000; // input=-2.763671875, output=-0.929433853419
			11'd1732: out = 32'b10000000000000000111011100100111; // input=-2.767578125, output=-0.930868121127
			11'd1733: out = 32'b10000000000000000111011101010101; // input=-2.771484375, output=-0.932288184932
			11'd1734: out = 32'b10000000000000000111011110000011; // input=-2.775390625, output=-0.933694023166
			11'd1735: out = 32'b10000000000000000111011110110001; // input=-2.779296875, output=-0.935085614378
			11'd1736: out = 32'b10000000000000000111011111011110; // input=-2.783203125, output=-0.936462937335
			11'd1737: out = 32'b10000000000000000111100000001011; // input=-2.787109375, output=-0.937825971019
			11'd1738: out = 32'b10000000000000000111100000110111; // input=-2.791015625, output=-0.939174694632
			11'd1739: out = 32'b10000000000000000111100001100011; // input=-2.794921875, output=-0.940509087596
			11'd1740: out = 32'b10000000000000000111100010001110; // input=-2.798828125, output=-0.941829129547
			11'd1741: out = 32'b10000000000000000111100010111001; // input=-2.802734375, output=-0.943134800345
			11'd1742: out = 32'b10000000000000000111100011100011; // input=-2.806640625, output=-0.944426080067
			11'd1743: out = 32'b10000000000000000111100100001101; // input=-2.810546875, output=-0.945702949008
			11'd1744: out = 32'b10000000000000000111100100110110; // input=-2.814453125, output=-0.946965387686
			11'd1745: out = 32'b10000000000000000111100101011111; // input=-2.818359375, output=-0.948213376837
			11'd1746: out = 32'b10000000000000000111100110000111; // input=-2.822265625, output=-0.949446897419
			11'd1747: out = 32'b10000000000000000111100110101111; // input=-2.826171875, output=-0.950665930609
			11'd1748: out = 32'b10000000000000000111100111010111; // input=-2.830078125, output=-0.951870457806
			11'd1749: out = 32'b10000000000000000111100111111110; // input=-2.833984375, output=-0.953060460632
			11'd1750: out = 32'b10000000000000000111101000100100; // input=-2.837890625, output=-0.954235920927
			11'd1751: out = 32'b10000000000000000111101001001010; // input=-2.841796875, output=-0.955396820757
			11'd1752: out = 32'b10000000000000000111101001110000; // input=-2.845703125, output=-0.956543142406
			11'd1753: out = 32'b10000000000000000111101010010101; // input=-2.849609375, output=-0.957674868384
			11'd1754: out = 32'b10000000000000000111101010111010; // input=-2.853515625, output=-0.958791981422
			11'd1755: out = 32'b10000000000000000111101011011110; // input=-2.857421875, output=-0.959894464473
			11'd1756: out = 32'b10000000000000000111101100000001; // input=-2.861328125, output=-0.960982300717
			11'd1757: out = 32'b10000000000000000111101100100101; // input=-2.865234375, output=-0.962055473552
			11'd1758: out = 32'b10000000000000000111101101000111; // input=-2.869140625, output=-0.963113966605
			11'd1759: out = 32'b10000000000000000111101101101010; // input=-2.873046875, output=-0.964157763723
			11'd1760: out = 32'b10000000000000000111101110001011; // input=-2.876953125, output=-0.965186848981
			11'd1761: out = 32'b10000000000000000111101110101100; // input=-2.880859375, output=-0.966201206674
			11'd1762: out = 32'b10000000000000000111101111001101; // input=-2.884765625, output=-0.967200821326
			11'd1763: out = 32'b10000000000000000111101111101110; // input=-2.888671875, output=-0.968185677683
			11'd1764: out = 32'b10000000000000000111110000001101; // input=-2.892578125, output=-0.969155760718
			11'd1765: out = 32'b10000000000000000111110000101101; // input=-2.896484375, output=-0.970111055629
			11'd1766: out = 32'b10000000000000000111110001001011; // input=-2.900390625, output=-0.971051547838
			11'd1767: out = 32'b10000000000000000111110001101010; // input=-2.904296875, output=-0.971977222996
			11'd1768: out = 32'b10000000000000000111110010001000; // input=-2.908203125, output=-0.972888066977
			11'd1769: out = 32'b10000000000000000111110010100101; // input=-2.912109375, output=-0.973784065883
			11'd1770: out = 32'b10000000000000000111110011000010; // input=-2.916015625, output=-0.974665206042
			11'd1771: out = 32'b10000000000000000111110011011110; // input=-2.919921875, output=-0.975531474009
			11'd1772: out = 32'b10000000000000000111110011111010; // input=-2.923828125, output=-0.976382856567
			11'd1773: out = 32'b10000000000000000111110100010110; // input=-2.927734375, output=-0.977219340723
			11'd1774: out = 32'b10000000000000000111110100110000; // input=-2.931640625, output=-0.978040913714
			11'd1775: out = 32'b10000000000000000111110101001011; // input=-2.935546875, output=-0.978847563005
			11'd1776: out = 32'b10000000000000000111110101100101; // input=-2.939453125, output=-0.979639276285
			11'd1777: out = 32'b10000000000000000111110101111110; // input=-2.943359375, output=-0.980416041476
			11'd1778: out = 32'b10000000000000000111110110010111; // input=-2.947265625, output=-0.981177846724
			11'd1779: out = 32'b10000000000000000111110110110000; // input=-2.951171875, output=-0.981924680406
			11'd1780: out = 32'b10000000000000000111110111001000; // input=-2.955078125, output=-0.982656531125
			11'd1781: out = 32'b10000000000000000111110111011111; // input=-2.958984375, output=-0.983373387714
			11'd1782: out = 32'b10000000000000000111110111110110; // input=-2.962890625, output=-0.984075239235
			11'd1783: out = 32'b10000000000000000111111000001101; // input=-2.966796875, output=-0.984762074979
			11'd1784: out = 32'b10000000000000000111111000100011; // input=-2.970703125, output=-0.985433884466
			11'd1785: out = 32'b10000000000000000111111000111000; // input=-2.974609375, output=-0.986090657443
			11'd1786: out = 32'b10000000000000000111111001001101; // input=-2.978515625, output=-0.986732383891
			11'd1787: out = 32'b10000000000000000111111001100010; // input=-2.982421875, output=-0.987359054016
			11'd1788: out = 32'b10000000000000000111111001110110; // input=-2.986328125, output=-0.987970658257
			11'd1789: out = 32'b10000000000000000111111010001001; // input=-2.990234375, output=-0.988567187281
			11'd1790: out = 32'b10000000000000000111111010011100; // input=-2.994140625, output=-0.989148631986
			11'd1791: out = 32'b10000000000000000111111010101111; // input=-2.998046875, output=-0.9897149835
			11'd1792: out = 32'b10000000000000000111111011000001; // input=-3.001953125, output=-0.990266233181
			11'd1793: out = 32'b10000000000000000111111011010011; // input=-3.005859375, output=-0.990802372617
			11'd1794: out = 32'b10000000000000000111111011100100; // input=-3.009765625, output=-0.991323393629
			11'd1795: out = 32'b10000000000000000111111011110100; // input=-3.013671875, output=-0.991829288265
			11'd1796: out = 32'b10000000000000000111111100000100; // input=-3.017578125, output=-0.992320048806
			11'd1797: out = 32'b10000000000000000111111100010100; // input=-3.021484375, output=-0.992795667765
			11'd1798: out = 32'b10000000000000000111111100100011; // input=-3.025390625, output=-0.993256137883
			11'd1799: out = 32'b10000000000000000111111100110010; // input=-3.029296875, output=-0.993701452134
			11'd1800: out = 32'b10000000000000000111111101000000; // input=-3.033203125, output=-0.994131603724
			11'd1801: out = 32'b10000000000000000111111101001101; // input=-3.037109375, output=-0.994546586089
			11'd1802: out = 32'b10000000000000000111111101011010; // input=-3.041015625, output=-0.994946392896
			11'd1803: out = 32'b10000000000000000111111101100111; // input=-3.044921875, output=-0.995331018046
			11'd1804: out = 32'b10000000000000000111111101110011; // input=-3.048828125, output=-0.995700455669
			11'd1805: out = 32'b10000000000000000111111101111111; // input=-3.052734375, output=-0.996054700128
			11'd1806: out = 32'b10000000000000000111111110001010; // input=-3.056640625, output=-0.996393746017
			11'd1807: out = 32'b10000000000000000111111110010100; // input=-3.060546875, output=-0.996717588164
			11'd1808: out = 32'b10000000000000000111111110011111; // input=-3.064453125, output=-0.997026221627
			11'd1809: out = 32'b10000000000000000111111110101000; // input=-3.068359375, output=-0.997319641697
			11'd1810: out = 32'b10000000000000000111111110110001; // input=-3.072265625, output=-0.997597843896
			11'd1811: out = 32'b10000000000000000111111110111010; // input=-3.076171875, output=-0.997860823979
			11'd1812: out = 32'b10000000000000000111111111000010; // input=-3.080078125, output=-0.998108577933
			11'd1813: out = 32'b10000000000000000111111111001010; // input=-3.083984375, output=-0.998341101979
			11'd1814: out = 32'b10000000000000000111111111010001; // input=-3.087890625, output=-0.998558392568
			11'd1815: out = 32'b10000000000000000111111111010111; // input=-3.091796875, output=-0.998760446384
			11'd1816: out = 32'b10000000000000000111111111011110; // input=-3.095703125, output=-0.998947260345
			11'd1817: out = 32'b10000000000000000111111111100011; // input=-3.099609375, output=-0.999118831599
			11'd1818: out = 32'b10000000000000000111111111101000; // input=-3.103515625, output=-0.99927515753
			11'd1819: out = 32'b10000000000000000111111111101101; // input=-3.107421875, output=-0.999416235751
			11'd1820: out = 32'b10000000000000000111111111110001; // input=-3.111328125, output=-0.99954206411
			11'd1821: out = 32'b10000000000000000111111111110101; // input=-3.115234375, output=-0.999652640687
			11'd1822: out = 32'b10000000000000000111111111111000; // input=-3.119140625, output=-0.999747963794
			11'd1823: out = 32'b10000000000000000111111111111010; // input=-3.123046875, output=-0.999828031977
			11'd1824: out = 32'b10000000000000000111111111111100; // input=-3.126953125, output=-0.999892844015
			11'd1825: out = 32'b10000000000000000111111111111110; // input=-3.130859375, output=-0.999942398918
			11'd1826: out = 32'b10000000000000000111111111111111; // input=-3.134765625, output=-0.999976695931
			11'd1827: out = 32'b10000000000000000111111111111111; // input=-3.138671875, output=-0.999995734529
			11'd1828: out = 32'b10000000000000000111111111111111; // input=-3.142578125, output=-0.999999514423
			11'd1829: out = 32'b10000000000000000111111111111111; // input=-3.146484375, output=-0.999988035555
			11'd1830: out = 32'b10000000000000000111111111111111; // input=-3.150390625, output=-0.999961298099
			11'd1831: out = 32'b10000000000000000111111111111101; // input=-3.154296875, output=-0.999919302465
			11'd1832: out = 32'b10000000000000000111111111111011; // input=-3.158203125, output=-0.999862049292
			11'd1833: out = 32'b10000000000000000111111111111001; // input=-3.162109375, output=-0.999789539454
			11'd1834: out = 32'b10000000000000000111111111110110; // input=-3.166015625, output=-0.999701774058
			11'd1835: out = 32'b10000000000000000111111111110011; // input=-3.169921875, output=-0.999598754443
			11'd1836: out = 32'b10000000000000000111111111101111; // input=-3.173828125, output=-0.999480482181
			11'd1837: out = 32'b10000000000000000111111111101011; // input=-3.177734375, output=-0.999346959076
			11'd1838: out = 32'b10000000000000000111111111100110; // input=-3.181640625, output=-0.999198187167
			11'd1839: out = 32'b10000000000000000111111111100000; // input=-3.185546875, output=-0.999034168722
			11'd1840: out = 32'b10000000000000000111111111011010; // input=-3.189453125, output=-0.998854906245
			11'd1841: out = 32'b10000000000000000111111111010100; // input=-3.193359375, output=-0.998660402471
			11'd1842: out = 32'b10000000000000000111111111001101; // input=-3.197265625, output=-0.998450660368
			11'd1843: out = 32'b10000000000000000111111111000110; // input=-3.201171875, output=-0.998225683137
			11'd1844: out = 32'b10000000000000000111111110111110; // input=-3.205078125, output=-0.997985474209
			11'd1845: out = 32'b10000000000000000111111110110110; // input=-3.208984375, output=-0.997730037251
			11'd1846: out = 32'b10000000000000000111111110101101; // input=-3.212890625, output=-0.997459376161
			11'd1847: out = 32'b10000000000000000111111110100011; // input=-3.216796875, output=-0.997173495067
			11'd1848: out = 32'b10000000000000000111111110011010; // input=-3.220703125, output=-0.996872398333
			11'd1849: out = 32'b10000000000000000111111110001111; // input=-3.224609375, output=-0.996556090553
			11'd1850: out = 32'b10000000000000000111111110000100; // input=-3.228515625, output=-0.996224576552
			11'd1851: out = 32'b10000000000000000111111101111001; // input=-3.232421875, output=-0.995877861391
			11'd1852: out = 32'b10000000000000000111111101101101; // input=-3.236328125, output=-0.995515950358
			11'd1853: out = 32'b10000000000000000111111101100001; // input=-3.240234375, output=-0.995138848977
			11'd1854: out = 32'b10000000000000000111111101010100; // input=-3.244140625, output=-0.994746563001
			11'd1855: out = 32'b10000000000000000111111101000111; // input=-3.248046875, output=-0.994339098417
			11'd1856: out = 32'b10000000000000000111111100111001; // input=-3.251953125, output=-0.993916461441
			11'd1857: out = 32'b10000000000000000111111100101010; // input=-3.255859375, output=-0.993478658524
			11'd1858: out = 32'b10000000000000000111111100011011; // input=-3.259765625, output=-0.993025696344
			11'd1859: out = 32'b10000000000000000111111100001100; // input=-3.263671875, output=-0.992557581813
			11'd1860: out = 32'b10000000000000000111111011111100; // input=-3.267578125, output=-0.992074322076
			11'd1861: out = 32'b10000000000000000111111011101100; // input=-3.271484375, output=-0.991575924504
			11'd1862: out = 32'b10000000000000000111111011011011; // input=-3.275390625, output=-0.991062396704
			11'd1863: out = 32'b10000000000000000111111011001010; // input=-3.279296875, output=-0.990533746511
			11'd1864: out = 32'b10000000000000000111111010111000; // input=-3.283203125, output=-0.989989981992
			11'd1865: out = 32'b10000000000000000111111010100110; // input=-3.287109375, output=-0.989431111444
			11'd1866: out = 32'b10000000000000000111111010010011; // input=-3.291015625, output=-0.988857143395
			11'd1867: out = 32'b10000000000000000111111010000000; // input=-3.294921875, output=-0.988268086602
			11'd1868: out = 32'b10000000000000000111111001101100; // input=-3.298828125, output=-0.987663950053
			11'd1869: out = 32'b10000000000000000111111001010111; // input=-3.302734375, output=-0.987044742969
			11'd1870: out = 32'b10000000000000000111111001000011; // input=-3.306640625, output=-0.986410474795
			11'd1871: out = 32'b10000000000000000111111000101101; // input=-3.310546875, output=-0.985761155212
			11'd1872: out = 32'b10000000000000000111111000011000; // input=-3.314453125, output=-0.985096794126
			11'd1873: out = 32'b10000000000000000111111000000001; // input=-3.318359375, output=-0.984417401675
			11'd1874: out = 32'b10000000000000000111110111101011; // input=-3.322265625, output=-0.983722988226
			11'd1875: out = 32'b10000000000000000111110111010011; // input=-3.326171875, output=-0.983013564374
			11'd1876: out = 32'b10000000000000000111110110111100; // input=-3.330078125, output=-0.982289140945
			11'd1877: out = 32'b10000000000000000111110110100011; // input=-3.333984375, output=-0.981549728992
			11'd1878: out = 32'b10000000000000000111110110001011; // input=-3.337890625, output=-0.980795339798
			11'd1879: out = 32'b10000000000000000111110101110001; // input=-3.341796875, output=-0.980025984873
			11'd1880: out = 32'b10000000000000000111110101011000; // input=-3.345703125, output=-0.979241675958
			11'd1881: out = 32'b10000000000000000111110100111110; // input=-3.349609375, output=-0.978442425019
			11'd1882: out = 32'b10000000000000000111110100100011; // input=-3.353515625, output=-0.977628244254
			11'd1883: out = 32'b10000000000000000111110100001000; // input=-3.357421875, output=-0.976799146083
			11'd1884: out = 32'b10000000000000000111110011101100; // input=-3.361328125, output=-0.97595514316
			11'd1885: out = 32'b10000000000000000111110011010000; // input=-3.365234375, output=-0.975096248362
			11'd1886: out = 32'b10000000000000000111110010110011; // input=-3.369140625, output=-0.974222474795
			11'd1887: out = 32'b10000000000000000111110010010110; // input=-3.373046875, output=-0.973333835791
			11'd1888: out = 32'b10000000000000000111110001111001; // input=-3.376953125, output=-0.972430344911
			11'd1889: out = 32'b10000000000000000111110001011011; // input=-3.380859375, output=-0.97151201594
			11'd1890: out = 32'b10000000000000000111110000111100; // input=-3.384765625, output=-0.970578862891
			11'd1891: out = 32'b10000000000000000111110000011101; // input=-3.388671875, output=-0.969630900003
			11'd1892: out = 32'b10000000000000000111101111111101; // input=-3.392578125, output=-0.96866814174
			11'd1893: out = 32'b10000000000000000111101111011101; // input=-3.396484375, output=-0.967690602793
			11'd1894: out = 32'b10000000000000000111101110111101; // input=-3.400390625, output=-0.966698298078
			11'd1895: out = 32'b10000000000000000111101110011100; // input=-3.404296875, output=-0.965691242737
			11'd1896: out = 32'b10000000000000000111101101111010; // input=-3.408203125, output=-0.964669452135
			11'd1897: out = 32'b10000000000000000111101101011000; // input=-3.412109375, output=-0.963632941864
			11'd1898: out = 32'b10000000000000000111101100110110; // input=-3.416015625, output=-0.96258172774
			11'd1899: out = 32'b10000000000000000111101100010011; // input=-3.419921875, output=-0.961515825803
			11'd1900: out = 32'b10000000000000000111101011110000; // input=-3.423828125, output=-0.960435252318
			11'd1901: out = 32'b10000000000000000111101011001100; // input=-3.427734375, output=-0.959340023773
			11'd1902: out = 32'b10000000000000000111101010100111; // input=-3.431640625, output=-0.958230156879
			11'd1903: out = 32'b10000000000000000111101010000010; // input=-3.435546875, output=-0.957105668571
			11'd1904: out = 32'b10000000000000000111101001011101; // input=-3.439453125, output=-0.955966576009
			11'd1905: out = 32'b10000000000000000111101000110111; // input=-3.443359375, output=-0.954812896573
			11'd1906: out = 32'b10000000000000000111101000010001; // input=-3.447265625, output=-0.953644647867
			11'd1907: out = 32'b10000000000000000111100111101010; // input=-3.451171875, output=-0.952461847717
			11'd1908: out = 32'b10000000000000000111100111000011; // input=-3.455078125, output=-0.951264514171
			11'd1909: out = 32'b10000000000000000111100110011011; // input=-3.458984375, output=-0.950052665499
			11'd1910: out = 32'b10000000000000000111100101110011; // input=-3.462890625, output=-0.948826320192
			11'd1911: out = 32'b10000000000000000111100101001010; // input=-3.466796875, output=-0.947585496963
			11'd1912: out = 32'b10000000000000000111100100100001; // input=-3.470703125, output=-0.946330214745
			11'd1913: out = 32'b10000000000000000111100011111000; // input=-3.474609375, output=-0.945060492692
			11'd1914: out = 32'b10000000000000000111100011001110; // input=-3.478515625, output=-0.943776350179
			11'd1915: out = 32'b10000000000000000111100010100011; // input=-3.482421875, output=-0.9424778068
			11'd1916: out = 32'b10000000000000000111100001111000; // input=-3.486328125, output=-0.94116488237
			11'd1917: out = 32'b10000000000000000111100001001101; // input=-3.490234375, output=-0.939837596921
			11'd1918: out = 32'b10000000000000000111100000100001; // input=-3.494140625, output=-0.938495970706
			11'd1919: out = 32'b10000000000000000111011111110100; // input=-3.498046875, output=-0.937140024198
			11'd1920: out = 32'b10000000000000000111011111000111; // input=-3.501953125, output=-0.935769778086
			11'd1921: out = 32'b10000000000000000111011110011010; // input=-3.505859375, output=-0.934385253279
			11'd1922: out = 32'b10000000000000000111011101101100; // input=-3.509765625, output=-0.932986470902
			11'd1923: out = 32'b10000000000000000111011100111110; // input=-3.513671875, output=-0.931573452299
			11'd1924: out = 32'b10000000000000000111011100001111; // input=-3.517578125, output=-0.930146219032
			11'd1925: out = 32'b10000000000000000111011011100000; // input=-3.521484375, output=-0.928704792878
			11'd1926: out = 32'b10000000000000000111011010110000; // input=-3.525390625, output=-0.927249195831
			11'd1927: out = 32'b10000000000000000111011010000000; // input=-3.529296875, output=-0.925779450103
			11'd1928: out = 32'b10000000000000000111011001001111; // input=-3.533203125, output=-0.924295578119
			11'd1929: out = 32'b10000000000000000111011000011110; // input=-3.537109375, output=-0.922797602521
			11'd1930: out = 32'b10000000000000000111010111101101; // input=-3.541015625, output=-0.921285546168
			11'd1931: out = 32'b10000000000000000111010110111011; // input=-3.544921875, output=-0.919759432131
			11'd1932: out = 32'b10000000000000000111010110001000; // input=-3.548828125, output=-0.918219283696
			11'd1933: out = 32'b10000000000000000111010101010101; // input=-3.552734375, output=-0.916665124365
			11'd1934: out = 32'b10000000000000000111010100100010; // input=-3.556640625, output=-0.915096977852
			11'd1935: out = 32'b10000000000000000111010011101110; // input=-3.560546875, output=-0.913514868085
			11'd1936: out = 32'b10000000000000000111010010111010; // input=-3.564453125, output=-0.911918819205
			11'd1937: out = 32'b10000000000000000111010010000101; // input=-3.568359375, output=-0.910308855566
			11'd1938: out = 32'b10000000000000000111010001010000; // input=-3.572265625, output=-0.908685001733
			11'd1939: out = 32'b10000000000000000111010000011010; // input=-3.576171875, output=-0.907047282486
			11'd1940: out = 32'b10000000000000000111001111100100; // input=-3.580078125, output=-0.905395722813
			11'd1941: out = 32'b10000000000000000111001110101101; // input=-3.583984375, output=-0.903730347915
			11'd1942: out = 32'b10000000000000000111001101110110; // input=-3.587890625, output=-0.902051183204
			11'd1943: out = 32'b10000000000000000111001100111111; // input=-3.591796875, output=-0.900358254301
			11'd1944: out = 32'b10000000000000000111001100000111; // input=-3.595703125, output=-0.89865158704
			11'd1945: out = 32'b10000000000000000111001011001111; // input=-3.599609375, output=-0.896931207461
			11'd1946: out = 32'b10000000000000000111001010010110; // input=-3.603515625, output=-0.895197141815
			11'd1947: out = 32'b10000000000000000111001001011101; // input=-3.607421875, output=-0.893449416562
			11'd1948: out = 32'b10000000000000000111001000100011; // input=-3.611328125, output=-0.89168805837
			11'd1949: out = 32'b10000000000000000111000111101001; // input=-3.615234375, output=-0.889913094116
			11'd1950: out = 32'b10000000000000000111000110101110; // input=-3.619140625, output=-0.888124550883
			11'd1951: out = 32'b10000000000000000111000101110011; // input=-3.623046875, output=-0.886322455962
			11'd1952: out = 32'b10000000000000000111000100111000; // input=-3.626953125, output=-0.88450683685
			11'd1953: out = 32'b10000000000000000111000011111100; // input=-3.630859375, output=-0.882677721253
			11'd1954: out = 32'b10000000000000000111000010111111; // input=-3.634765625, output=-0.880835137079
			11'd1955: out = 32'b10000000000000000111000010000010; // input=-3.638671875, output=-0.878979112445
			11'd1956: out = 32'b10000000000000000111000001000101; // input=-3.642578125, output=-0.877109675671
			11'd1957: out = 32'b10000000000000000111000000000111; // input=-3.646484375, output=-0.875226855283
			11'd1958: out = 32'b10000000000000000110111111001001; // input=-3.650390625, output=-0.87333068001
			11'd1959: out = 32'b10000000000000000110111110001011; // input=-3.654296875, output=-0.871421178785
			11'd1960: out = 32'b10000000000000000110111101001100; // input=-3.658203125, output=-0.869498380745
			11'd1961: out = 32'b10000000000000000110111100001100; // input=-3.662109375, output=-0.867562315229
			11'd1962: out = 32'b10000000000000000110111011001100; // input=-3.666015625, output=-0.86561301178
			11'd1963: out = 32'b10000000000000000110111010001100; // input=-3.669921875, output=-0.863650500142
			11'd1964: out = 32'b10000000000000000110111001001011; // input=-3.673828125, output=-0.861674810259
			11'd1965: out = 32'b10000000000000000110111000001010; // input=-3.677734375, output=-0.859685972279
			11'd1966: out = 32'b10000000000000000110110111001001; // input=-3.681640625, output=-0.857684016548
			11'd1967: out = 32'b10000000000000000110110110000111; // input=-3.685546875, output=-0.855668973615
			11'd1968: out = 32'b10000000000000000110110101000100; // input=-3.689453125, output=-0.853640874226
			11'd1969: out = 32'b10000000000000000110110100000001; // input=-3.693359375, output=-0.851599749328
			11'd1970: out = 32'b10000000000000000110110010111110; // input=-3.697265625, output=-0.849545630065
			11'd1971: out = 32'b10000000000000000110110001111010; // input=-3.701171875, output=-0.847478547781
			11'd1972: out = 32'b10000000000000000110110000110110; // input=-3.705078125, output=-0.845398534017
			11'd1973: out = 32'b10000000000000000110101111110001; // input=-3.708984375, output=-0.843305620512
			11'd1974: out = 32'b10000000000000000110101110101100; // input=-3.712890625, output=-0.8411998392
			11'd1975: out = 32'b10000000000000000110101101100111; // input=-3.716796875, output=-0.839081222214
			11'd1976: out = 32'b10000000000000000110101100100001; // input=-3.720703125, output=-0.83694980188
			11'd1977: out = 32'b10000000000000000110101011011011; // input=-3.724609375, output=-0.834805610723
			11'd1978: out = 32'b10000000000000000110101010010100; // input=-3.728515625, output=-0.832648681459
			11'd1979: out = 32'b10000000000000000110101001001101; // input=-3.732421875, output=-0.830479047
			11'd1980: out = 32'b10000000000000000110101000000110; // input=-3.736328125, output=-0.828296740453
			11'd1981: out = 32'b10000000000000000110100110111110; // input=-3.740234375, output=-0.826101795117
			11'd1982: out = 32'b10000000000000000110100101110101; // input=-3.744140625, output=-0.823894244484
			11'd1983: out = 32'b10000000000000000110100100101101; // input=-3.748046875, output=-0.821674122238
			11'd1984: out = 32'b10000000000000000110100011100011; // input=-3.751953125, output=-0.819441462256
			11'd1985: out = 32'b10000000000000000110100010011010; // input=-3.755859375, output=-0.817196298606
			11'd1986: out = 32'b10000000000000000110100001010000; // input=-3.759765625, output=-0.814938665546
			11'd1987: out = 32'b10000000000000000110100000000110; // input=-3.763671875, output=-0.812668597524
			11'd1988: out = 32'b10000000000000000110011110111011; // input=-3.767578125, output=-0.810386129179
			11'd1989: out = 32'b10000000000000000110011101110000; // input=-3.771484375, output=-0.808091295339
			11'd1990: out = 32'b10000000000000000110011100100100; // input=-3.775390625, output=-0.80578413102
			11'd1991: out = 32'b10000000000000000110011011011000; // input=-3.779296875, output=-0.803464671426
			11'd1992: out = 32'b10000000000000000110011010001100; // input=-3.783203125, output=-0.801132951951
			11'd1993: out = 32'b10000000000000000110011000111111; // input=-3.787109375, output=-0.798789008172
			11'd1994: out = 32'b10000000000000000110010111110010; // input=-3.791015625, output=-0.796432875855
			11'd1995: out = 32'b10000000000000000110010110100100; // input=-3.794921875, output=-0.794064590953
			11'd1996: out = 32'b10000000000000000110010101010110; // input=-3.798828125, output=-0.791684189602
			11'd1997: out = 32'b10000000000000000110010100001000; // input=-3.802734375, output=-0.789291708124
			11'd1998: out = 32'b10000000000000000110010010111001; // input=-3.806640625, output=-0.786887183026
			11'd1999: out = 32'b10000000000000000110010001101010; // input=-3.810546875, output=-0.784470650998
			11'd2000: out = 32'b10000000000000000110010000011010; // input=-3.814453125, output=-0.782042148913
			11'd2001: out = 32'b10000000000000000110001111001010; // input=-3.818359375, output=-0.779601713826
			11'd2002: out = 32'b10000000000000000110001101111010; // input=-3.822265625, output=-0.777149382977
			11'd2003: out = 32'b10000000000000000110001100101001; // input=-3.826171875, output=-0.774685193784
			11'd2004: out = 32'b10000000000000000110001011011000; // input=-3.830078125, output=-0.772209183849
			11'd2005: out = 32'b10000000000000000110001010000110; // input=-3.833984375, output=-0.769721390951
			11'd2006: out = 32'b10000000000000000110001000110100; // input=-3.837890625, output=-0.767221853052
			11'd2007: out = 32'b10000000000000000110000111100010; // input=-3.841796875, output=-0.764710608291
			11'd2008: out = 32'b10000000000000000110000110001111; // input=-3.845703125, output=-0.762187694988
			11'd2009: out = 32'b10000000000000000110000100111100; // input=-3.849609375, output=-0.759653151638
			11'd2010: out = 32'b10000000000000000110000011101001; // input=-3.853515625, output=-0.757107016915
			11'd2011: out = 32'b10000000000000000110000010010101; // input=-3.857421875, output=-0.754549329671
			11'd2012: out = 32'b10000000000000000110000001000001; // input=-3.861328125, output=-0.751980128932
			11'd2013: out = 32'b10000000000000000101111111101100; // input=-3.865234375, output=-0.749399453902
			11'd2014: out = 32'b10000000000000000101111110010111; // input=-3.869140625, output=-0.746807343958
			11'd2015: out = 32'b10000000000000000101111101000010; // input=-3.873046875, output=-0.744203838653
			11'd2016: out = 32'b10000000000000000101111011101100; // input=-3.876953125, output=-0.741588977713
			11'd2017: out = 32'b10000000000000000101111010010110; // input=-3.880859375, output=-0.738962801038
			11'd2018: out = 32'b10000000000000000101111001000000; // input=-3.884765625, output=-0.736325348699
			11'd2019: out = 32'b10000000000000000101110111101001; // input=-3.888671875, output=-0.733676660942
			11'd2020: out = 32'b10000000000000000101110110010010; // input=-3.892578125, output=-0.731016778181
			11'd2021: out = 32'b10000000000000000101110100111010; // input=-3.896484375, output=-0.728345741004
			11'd2022: out = 32'b10000000000000000101110011100011; // input=-3.900390625, output=-0.725663590167
			11'd2023: out = 32'b10000000000000000101110010001010; // input=-3.904296875, output=-0.722970366596
			11'd2024: out = 32'b10000000000000000101110000110010; // input=-3.908203125, output=-0.720266111387
			11'd2025: out = 32'b10000000000000000101101111011001; // input=-3.912109375, output=-0.717550865803
			11'd2026: out = 32'b10000000000000000101101101111111; // input=-3.916015625, output=-0.714824671276
			11'd2027: out = 32'b10000000000000000101101100100110; // input=-3.919921875, output=-0.712087569404
			11'd2028: out = 32'b10000000000000000101101011001100; // input=-3.923828125, output=-0.709339601952
			11'd2029: out = 32'b10000000000000000101101001110001; // input=-3.927734375, output=-0.70658081085
			11'd2030: out = 32'b10000000000000000101101000010110; // input=-3.931640625, output=-0.703811238194
			11'd2031: out = 32'b10000000000000000101100110111011; // input=-3.935546875, output=-0.701030926245
			11'd2032: out = 32'b10000000000000000101100101100000; // input=-3.939453125, output=-0.698239917426
			11'd2033: out = 32'b10000000000000000101100100000100; // input=-3.943359375, output=-0.695438254325
			11'd2034: out = 32'b10000000000000000101100010101000; // input=-3.947265625, output=-0.692625979692
			11'd2035: out = 32'b10000000000000000101100001001011; // input=-3.951171875, output=-0.689803136439
			11'd2036: out = 32'b10000000000000000101011111101111; // input=-3.955078125, output=-0.686969767639
			11'd2037: out = 32'b10000000000000000101011110010001; // input=-3.958984375, output=-0.684125916525
			11'd2038: out = 32'b10000000000000000101011100110100; // input=-3.962890625, output=-0.681271626491
			11'd2039: out = 32'b10000000000000000101011011010110; // input=-3.966796875, output=-0.678406941091
			11'd2040: out = 32'b10000000000000000101011001111000; // input=-3.970703125, output=-0.675531904035
			11'd2041: out = 32'b10000000000000000101011000011001; // input=-3.974609375, output=-0.672646559194
			11'd2042: out = 32'b10000000000000000101010110111010; // input=-3.978515625, output=-0.669750950593
			11'd2043: out = 32'b10000000000000000101010101011011; // input=-3.982421875, output=-0.666845122418
			11'd2044: out = 32'b10000000000000000101010011111100; // input=-3.986328125, output=-0.663929119006
			11'd2045: out = 32'b10000000000000000101010010011100; // input=-3.990234375, output=-0.661002984852
			11'd2046: out = 32'b10000000000000000101010000111100; // input=-3.994140625, output=-0.658066764607
			11'd2047: out = 32'b10000000000000000101001111011011; // input=-3.998046875, output=-0.655120503072
		endcase
	end
	converter U0 (a, index);

endmodule