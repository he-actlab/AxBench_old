// Developed by: 	Amir Yazdanbakhsh
// Email: 			a.yazdanbakhsh@gatech.edu
// Date:			December 5, 2014

`timescale 1ns / 1ps

module gaussian_rom(addr, data_out);
	
	input  		[4:0]  addr;
	output reg 	[15:0] data_out;

	always @(addr)
	begin
		case(addr)
			5'd0: 		data_out <= 16'b0000_0000_0011_0100; // 2/159
			5'd1: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd2: 		data_out <= 16'b0000_0000_1000_0001; // 5/159
			5'd3: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd4: 		data_out <= 16'b0000_0000_0011_0100; // 2/159
			5'd5: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd6: 		data_out <= 16'b0000_0000_1110_1000; // 9/159
			5'd7: 		data_out <= 16'b0000_0001_0011_0101; // 12/159
			5'd8: 		data_out <= 16'b0000_0000_1110_1000; // 9/159
			5'd9:   	data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd10: 		data_out <= 16'b0000_0000_1000_0001; // 5/159
			5'd11: 		data_out <= 16'b0000_0001_0011_0101; // 12/159
			5'd12: 		data_out <= 16'b0000_0001_1000_0010; // 15/159
			5'd13: 		data_out <= 16'b0000_0001_0011_0101; // 12/159
			5'd14: 		data_out <= 16'b0000_0000_1000_0001; // 5/159
			5'd15: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd16: 		data_out <= 16'b0000_0000_1110_1000; // 9/159
			5'd17: 		data_out <= 16'b0000_0001_0011_0101; // 12/159
			5'd18: 		data_out <= 16'b0000_0000_1110_1000; // 9/159
			5'd19: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd20: 		data_out <= 16'b0000_0000_0011_0100; // 2/159
			5'd21: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd22: 		data_out <= 16'b0000_0000_1000_0001; // 5/159
			5'd23: 		data_out <= 16'b0000_0000_0110_0111; // 4/159
			5'd24: 		data_out <= 16'b0000_0000_0011_0100; // 2/159
			default: 	data_out <= 16'b0000_0000_0000_0000;
		endcase
	end
	
endmodule