// Developed by: Amir Yazdanbakhsh
// Email: a.yazdanbakhsh@gatech.edu

`timescale 1ns/1ps
module acos_lut(a, out);
	input  [31:0] a;
	output reg [31:0] out;
	wire   [10:0] index;

	always @(index)
	begin
		case(index)
			11'd0: out = 32'b00000000000000001100100100000000; // input=0.00048828125, output=1.57030804553
			11'd1: out = 32'b00000000000000001100100011100000; // input=0.00146484375, output=1.56933148252
			11'd2: out = 32'b00000000000000001100100011000000; // input=0.00244140625, output=1.56835491812
			11'd3: out = 32'b00000000000000001100100010100000; // input=0.00341796875, output=1.56737835139
			11'd4: out = 32'b00000000000000001100100010000000; // input=0.00439453125, output=1.5664017814
			11'd5: out = 32'b00000000000000001100100001100000; // input=0.00537109375, output=1.56542520722
			11'd6: out = 32'b00000000000000001100100001000000; // input=0.00634765625, output=1.56444862792
			11'd7: out = 32'b00000000000000001100100000100000; // input=0.00732421875, output=1.56347204256
			11'd8: out = 32'b00000000000000001100100000000000; // input=0.00830078125, output=1.56249545022
			11'd9: out = 32'b00000000000000001100011111100000; // input=0.00927734375, output=1.56151884996
			11'd10: out = 32'b00000000000000001100011111000000; // input=0.01025390625, output=1.56054224085
			11'd11: out = 32'b00000000000000001100011110100000; // input=0.01123046875, output=1.55956562196
			11'd12: out = 32'b00000000000000001100011110000000; // input=0.01220703125, output=1.55858899236
			11'd13: out = 32'b00000000000000001100011101100000; // input=0.01318359375, output=1.55761235111
			11'd14: out = 32'b00000000000000001100011101000000; // input=0.01416015625, output=1.55663569729
			11'd15: out = 32'b00000000000000001100011100100000; // input=0.01513671875, output=1.55565902996
			11'd16: out = 32'b00000000000000001100011100000000; // input=0.01611328125, output=1.55468234819
			11'd17: out = 32'b00000000000000001100011011100000; // input=0.01708984375, output=1.55370565105
			11'd18: out = 32'b00000000000000001100011011000000; // input=0.01806640625, output=1.5527289376
			11'd19: out = 32'b00000000000000001100011010100000; // input=0.01904296875, output=1.55175220692
			11'd20: out = 32'b00000000000000001100011010000000; // input=0.02001953125, output=1.55077545806
			11'd21: out = 32'b00000000000000001100011001100000; // input=0.02099609375, output=1.5497986901
			11'd22: out = 32'b00000000000000001100011001000000; // input=0.02197265625, output=1.5488219021
			11'd23: out = 32'b00000000000000001100011000100000; // input=0.02294921875, output=1.54784509314
			11'd24: out = 32'b00000000000000001100011000000000; // input=0.02392578125, output=1.54686826227
			11'd25: out = 32'b00000000000000001100010111100000; // input=0.02490234375, output=1.54589140856
			11'd26: out = 32'b00000000000000001100010111000000; // input=0.02587890625, output=1.54491453108
			11'd27: out = 32'b00000000000000001100010110100000; // input=0.02685546875, output=1.5439376289
			11'd28: out = 32'b00000000000000001100010110000000; // input=0.02783203125, output=1.54296070107
			11'd29: out = 32'b00000000000000001100010101100000; // input=0.02880859375, output=1.54198374668
			11'd30: out = 32'b00000000000000001100010101000000; // input=0.02978515625, output=1.54100676477
			11'd31: out = 32'b00000000000000001100010100100000; // input=0.03076171875, output=1.54002975443
			11'd32: out = 32'b00000000000000001100010100000000; // input=0.03173828125, output=1.5390527147
			11'd33: out = 32'b00000000000000001100010011100000; // input=0.03271484375, output=1.53807564466
			11'd34: out = 32'b00000000000000001100010011000000; // input=0.03369140625, output=1.53709854337
			11'd35: out = 32'b00000000000000001100010010100000; // input=0.03466796875, output=1.5361214099
			11'd36: out = 32'b00000000000000001100010010000000; // input=0.03564453125, output=1.5351442433
			11'd37: out = 32'b00000000000000001100010001100000; // input=0.03662109375, output=1.53416704265
			11'd38: out = 32'b00000000000000001100010001000000; // input=0.03759765625, output=1.533189807
			11'd39: out = 32'b00000000000000001100010000100000; // input=0.03857421875, output=1.53221253542
			11'd40: out = 32'b00000000000000001100010000000000; // input=0.03955078125, output=1.53123522697
			11'd41: out = 32'b00000000000000001100001111011111; // input=0.04052734375, output=1.53025788071
			11'd42: out = 32'b00000000000000001100001110111111; // input=0.04150390625, output=1.52928049571
			11'd43: out = 32'b00000000000000001100001110011111; // input=0.04248046875, output=1.52830307102
			11'd44: out = 32'b00000000000000001100001101111111; // input=0.04345703125, output=1.52732560571
			11'd45: out = 32'b00000000000000001100001101011111; // input=0.04443359375, output=1.52634809884
			11'd46: out = 32'b00000000000000001100001100111111; // input=0.04541015625, output=1.52537054947
			11'd47: out = 32'b00000000000000001100001100011111; // input=0.04638671875, output=1.52439295665
			11'd48: out = 32'b00000000000000001100001011111111; // input=0.04736328125, output=1.52341531946
			11'd49: out = 32'b00000000000000001100001011011111; // input=0.04833984375, output=1.52243763694
			11'd50: out = 32'b00000000000000001100001010111111; // input=0.04931640625, output=1.52145990816
			11'd51: out = 32'b00000000000000001100001010011111; // input=0.05029296875, output=1.52048213218
			11'd52: out = 32'b00000000000000001100001001111111; // input=0.05126953125, output=1.51950430805
			11'd53: out = 32'b00000000000000001100001001011111; // input=0.05224609375, output=1.51852643484
			11'd54: out = 32'b00000000000000001100001000111111; // input=0.05322265625, output=1.51754851159
			11'd55: out = 32'b00000000000000001100001000011111; // input=0.05419921875, output=1.51657053737
			11'd56: out = 32'b00000000000000001100000111111111; // input=0.05517578125, output=1.51559251124
			11'd57: out = 32'b00000000000000001100000111011111; // input=0.05615234375, output=1.51461443224
			11'd58: out = 32'b00000000000000001100000110111111; // input=0.05712890625, output=1.51363629943
			11'd59: out = 32'b00000000000000001100000110011111; // input=0.05810546875, output=1.51265811188
			11'd60: out = 32'b00000000000000001100000101111111; // input=0.05908203125, output=1.51167986863
			11'd61: out = 32'b00000000000000001100000101011111; // input=0.06005859375, output=1.51070156874
			11'd62: out = 32'b00000000000000001100000100111111; // input=0.06103515625, output=1.50972321126
			11'd63: out = 32'b00000000000000001100000100011111; // input=0.06201171875, output=1.50874479525
			11'd64: out = 32'b00000000000000001100000011111110; // input=0.06298828125, output=1.50776631976
			11'd65: out = 32'b00000000000000001100000011011110; // input=0.06396484375, output=1.50678778383
			11'd66: out = 32'b00000000000000001100000010111110; // input=0.06494140625, output=1.50580918653
			11'd67: out = 32'b00000000000000001100000010011110; // input=0.06591796875, output=1.5048305269
			11'd68: out = 32'b00000000000000001100000001111110; // input=0.06689453125, output=1.503851804
			11'd69: out = 32'b00000000000000001100000001011110; // input=0.06787109375, output=1.50287301687
			11'd70: out = 32'b00000000000000001100000000111110; // input=0.06884765625, output=1.50189416456
			11'd71: out = 32'b00000000000000001100000000011110; // input=0.06982421875, output=1.50091524612
			11'd72: out = 32'b00000000000000001011111111111110; // input=0.07080078125, output=1.49993626061
			11'd73: out = 32'b00000000000000001011111111011110; // input=0.07177734375, output=1.49895720706
			11'd74: out = 32'b00000000000000001011111110111110; // input=0.07275390625, output=1.49797808453
			11'd75: out = 32'b00000000000000001011111110011110; // input=0.07373046875, output=1.49699889206
			11'd76: out = 32'b00000000000000001011111101111110; // input=0.07470703125, output=1.49601962869
			11'd77: out = 32'b00000000000000001011111101011101; // input=0.07568359375, output=1.49504029348
			11'd78: out = 32'b00000000000000001011111100111101; // input=0.07666015625, output=1.49406088547
			11'd79: out = 32'b00000000000000001011111100011101; // input=0.07763671875, output=1.4930814037
			11'd80: out = 32'b00000000000000001011111011111101; // input=0.07861328125, output=1.49210184722
			11'd81: out = 32'b00000000000000001011111011011101; // input=0.07958984375, output=1.49112221506
			11'd82: out = 32'b00000000000000001011111010111101; // input=0.08056640625, output=1.49014250628
			11'd83: out = 32'b00000000000000001011111010011101; // input=0.08154296875, output=1.4891627199
			11'd84: out = 32'b00000000000000001011111001111101; // input=0.08251953125, output=1.48818285498
			11'd85: out = 32'b00000000000000001011111001011101; // input=0.08349609375, output=1.48720291055
			11'd86: out = 32'b00000000000000001011111000111101; // input=0.08447265625, output=1.48622288565
			11'd87: out = 32'b00000000000000001011111000011100; // input=0.08544921875, output=1.48524277933
			11'd88: out = 32'b00000000000000001011110111111100; // input=0.08642578125, output=1.48426259061
			11'd89: out = 32'b00000000000000001011110111011100; // input=0.08740234375, output=1.48328231853
			11'd90: out = 32'b00000000000000001011110110111100; // input=0.08837890625, output=1.48230196214
			11'd91: out = 32'b00000000000000001011110110011100; // input=0.08935546875, output=1.48132152047
			11'd92: out = 32'b00000000000000001011110101111100; // input=0.09033203125, output=1.48034099255
			11'd93: out = 32'b00000000000000001011110101011100; // input=0.09130859375, output=1.47936037742
			11'd94: out = 32'b00000000000000001011110100111100; // input=0.09228515625, output=1.47837967411
			11'd95: out = 32'b00000000000000001011110100011011; // input=0.09326171875, output=1.47739888165
			11'd96: out = 32'b00000000000000001011110011111011; // input=0.09423828125, output=1.47641799908
			11'd97: out = 32'b00000000000000001011110011011011; // input=0.09521484375, output=1.47543702542
			11'd98: out = 32'b00000000000000001011110010111011; // input=0.09619140625, output=1.47445595971
			11'd99: out = 32'b00000000000000001011110010011011; // input=0.09716796875, output=1.47347480098
			11'd100: out = 32'b00000000000000001011110001111011; // input=0.09814453125, output=1.47249354825
			11'd101: out = 32'b00000000000000001011110001011011; // input=0.09912109375, output=1.47151220056
			11'd102: out = 32'b00000000000000001011110000111010; // input=0.10009765625, output=1.47053075692
			11'd103: out = 32'b00000000000000001011110000011010; // input=0.10107421875, output=1.46954921638
			11'd104: out = 32'b00000000000000001011101111111010; // input=0.10205078125, output=1.46856757794
			11'd105: out = 32'b00000000000000001011101111011010; // input=0.10302734375, output=1.46758584064
			11'd106: out = 32'b00000000000000001011101110111010; // input=0.10400390625, output=1.4666040035
			11'd107: out = 32'b00000000000000001011101110011010; // input=0.10498046875, output=1.46562206555
			11'd108: out = 32'b00000000000000001011101101111001; // input=0.10595703125, output=1.4646400258
			11'd109: out = 32'b00000000000000001011101101011001; // input=0.10693359375, output=1.46365788327
			11'd110: out = 32'b00000000000000001011101100111001; // input=0.10791015625, output=1.46267563699
			11'd111: out = 32'b00000000000000001011101100011001; // input=0.10888671875, output=1.46169328597
			11'd112: out = 32'b00000000000000001011101011111001; // input=0.10986328125, output=1.46071082924
			11'd113: out = 32'b00000000000000001011101011011000; // input=0.11083984375, output=1.45972826581
			11'd114: out = 32'b00000000000000001011101010111000; // input=0.11181640625, output=1.45874559469
			11'd115: out = 32'b00000000000000001011101010011000; // input=0.11279296875, output=1.45776281491
			11'd116: out = 32'b00000000000000001011101001111000; // input=0.11376953125, output=1.45677992547
			11'd117: out = 32'b00000000000000001011101001011000; // input=0.11474609375, output=1.45579692539
			11'd118: out = 32'b00000000000000001011101000110111; // input=0.11572265625, output=1.45481381369
			11'd119: out = 32'b00000000000000001011101000010111; // input=0.11669921875, output=1.45383058936
			11'd120: out = 32'b00000000000000001011100111110111; // input=0.11767578125, output=1.45284725144
			11'd121: out = 32'b00000000000000001011100111010111; // input=0.11865234375, output=1.45186379891
			11'd122: out = 32'b00000000000000001011100110110110; // input=0.11962890625, output=1.4508802308
			11'd123: out = 32'b00000000000000001011100110010110; // input=0.12060546875, output=1.4498965461
			11'd124: out = 32'b00000000000000001011100101110110; // input=0.12158203125, output=1.44891274383
			11'd125: out = 32'b00000000000000001011100101010110; // input=0.12255859375, output=1.447928823
			11'd126: out = 32'b00000000000000001011100100110101; // input=0.12353515625, output=1.4469447826
			11'd127: out = 32'b00000000000000001011100100010101; // input=0.12451171875, output=1.44596062163
			11'd128: out = 32'b00000000000000001011100011110101; // input=0.12548828125, output=1.44497633911
			11'd129: out = 32'b00000000000000001011100011010101; // input=0.12646484375, output=1.44399193403
			11'd130: out = 32'b00000000000000001011100010110100; // input=0.12744140625, output=1.44300740539
			11'd131: out = 32'b00000000000000001011100010010100; // input=0.12841796875, output=1.44202275218
			11'd132: out = 32'b00000000000000001011100001110100; // input=0.12939453125, output=1.44103797342
			11'd133: out = 32'b00000000000000001011100001010100; // input=0.13037109375, output=1.44005306809
			11'd134: out = 32'b00000000000000001011100000110011; // input=0.13134765625, output=1.4390680352
			11'd135: out = 32'b00000000000000001011100000010011; // input=0.13232421875, output=1.43808287372
			11'd136: out = 32'b00000000000000001011011111110011; // input=0.13330078125, output=1.43709758266
			11'd137: out = 32'b00000000000000001011011111010011; // input=0.13427734375, output=1.43611216102
			11'd138: out = 32'b00000000000000001011011110110010; // input=0.13525390625, output=1.43512660777
			11'd139: out = 32'b00000000000000001011011110010010; // input=0.13623046875, output=1.43414092191
			11'd140: out = 32'b00000000000000001011011101110010; // input=0.13720703125, output=1.43315510243
			11'd141: out = 32'b00000000000000001011011101010001; // input=0.13818359375, output=1.43216914831
			11'd142: out = 32'b00000000000000001011011100110001; // input=0.13916015625, output=1.43118305855
			11'd143: out = 32'b00000000000000001011011100010001; // input=0.14013671875, output=1.43019683212
			11'd144: out = 32'b00000000000000001011011011110000; // input=0.14111328125, output=1.42921046801
			11'd145: out = 32'b00000000000000001011011011010000; // input=0.14208984375, output=1.4282239652
			11'd146: out = 32'b00000000000000001011011010110000; // input=0.14306640625, output=1.42723732268
			11'd147: out = 32'b00000000000000001011011010001111; // input=0.14404296875, output=1.42625053942
			11'd148: out = 32'b00000000000000001011011001101111; // input=0.14501953125, output=1.42526361439
			11'd149: out = 32'b00000000000000001011011001001111; // input=0.14599609375, output=1.42427654659
			11'd150: out = 32'b00000000000000001011011000101110; // input=0.14697265625, output=1.42328933498
			11'd151: out = 32'b00000000000000001011011000001110; // input=0.14794921875, output=1.42230197854
			11'd152: out = 32'b00000000000000001011010111101110; // input=0.14892578125, output=1.42131447624
			11'd153: out = 32'b00000000000000001011010111001101; // input=0.14990234375, output=1.42032682706
			11'd154: out = 32'b00000000000000001011010110101101; // input=0.15087890625, output=1.41933902995
			11'd155: out = 32'b00000000000000001011010110001101; // input=0.15185546875, output=1.41835108391
			11'd156: out = 32'b00000000000000001011010101101100; // input=0.15283203125, output=1.41736298788
			11'd157: out = 32'b00000000000000001011010101001100; // input=0.15380859375, output=1.41637474084
			11'd158: out = 32'b00000000000000001011010100101011; // input=0.15478515625, output=1.41538634176
			11'd159: out = 32'b00000000000000001011010100001011; // input=0.15576171875, output=1.41439778959
			11'd160: out = 32'b00000000000000001011010011101011; // input=0.15673828125, output=1.4134090833
			11'd161: out = 32'b00000000000000001011010011001010; // input=0.15771484375, output=1.41242022185
			11'd162: out = 32'b00000000000000001011010010101010; // input=0.15869140625, output=1.4114312042
			11'd163: out = 32'b00000000000000001011010010001001; // input=0.15966796875, output=1.41044202931
			11'd164: out = 32'b00000000000000001011010001101001; // input=0.16064453125, output=1.40945269613
			11'd165: out = 32'b00000000000000001011010001001001; // input=0.16162109375, output=1.40846320363
			11'd166: out = 32'b00000000000000001011010000101000; // input=0.16259765625, output=1.40747355074
			11'd167: out = 32'b00000000000000001011010000001000; // input=0.16357421875, output=1.40648373644
			11'd168: out = 32'b00000000000000001011001111100111; // input=0.16455078125, output=1.40549375965
			11'd169: out = 32'b00000000000000001011001111000111; // input=0.16552734375, output=1.40450361935
			11'd170: out = 32'b00000000000000001011001110100110; // input=0.16650390625, output=1.40351331446
			11'd171: out = 32'b00000000000000001011001110000110; // input=0.16748046875, output=1.40252284395
			11'd172: out = 32'b00000000000000001011001101100101; // input=0.16845703125, output=1.40153220675
			11'd173: out = 32'b00000000000000001011001101000101; // input=0.16943359375, output=1.40054140181
			11'd174: out = 32'b00000000000000001011001100100100; // input=0.17041015625, output=1.39955042807
			11'd175: out = 32'b00000000000000001011001100000100; // input=0.17138671875, output=1.39855928446
			11'd176: out = 32'b00000000000000001011001011100100; // input=0.17236328125, output=1.39756796994
			11'd177: out = 32'b00000000000000001011001011000011; // input=0.17333984375, output=1.39657648342
			11'd178: out = 32'b00000000000000001011001010100011; // input=0.17431640625, output=1.39558482386
			11'd179: out = 32'b00000000000000001011001010000010; // input=0.17529296875, output=1.39459299018
			11'd180: out = 32'b00000000000000001011001001100010; // input=0.17626953125, output=1.39360098132
			11'd181: out = 32'b00000000000000001011001001000001; // input=0.17724609375, output=1.3926087962
			11'd182: out = 32'b00000000000000001011001000100000; // input=0.17822265625, output=1.39161643376
			11'd183: out = 32'b00000000000000001011001000000000; // input=0.17919921875, output=1.39062389291
			11'd184: out = 32'b00000000000000001011000111011111; // input=0.18017578125, output=1.3896311726
			11'd185: out = 32'b00000000000000001011000110111111; // input=0.18115234375, output=1.38863827173
			11'd186: out = 32'b00000000000000001011000110011110; // input=0.18212890625, output=1.38764518924
			11'd187: out = 32'b00000000000000001011000101111110; // input=0.18310546875, output=1.38665192404
			11'd188: out = 32'b00000000000000001011000101011101; // input=0.18408203125, output=1.38565847506
			11'd189: out = 32'b00000000000000001011000100111101; // input=0.18505859375, output=1.3846648412
			11'd190: out = 32'b00000000000000001011000100011100; // input=0.18603515625, output=1.38367102139
			11'd191: out = 32'b00000000000000001011000011111100; // input=0.18701171875, output=1.38267701453
			11'd192: out = 32'b00000000000000001011000011011011; // input=0.18798828125, output=1.38168281954
			11'd193: out = 32'b00000000000000001011000010111010; // input=0.18896484375, output=1.38068843533
			11'd194: out = 32'b00000000000000001011000010011010; // input=0.18994140625, output=1.37969386081
			11'd195: out = 32'b00000000000000001011000001111001; // input=0.19091796875, output=1.37869909488
			11'd196: out = 32'b00000000000000001011000001011001; // input=0.19189453125, output=1.37770413645
			11'd197: out = 32'b00000000000000001011000000111000; // input=0.19287109375, output=1.37670898442
			11'd198: out = 32'b00000000000000001011000000010111; // input=0.19384765625, output=1.37571363769
			11'd199: out = 32'b00000000000000001010111111110111; // input=0.19482421875, output=1.37471809517
			11'd200: out = 32'b00000000000000001010111111010110; // input=0.19580078125, output=1.37372235573
			11'd201: out = 32'b00000000000000001010111110110101; // input=0.19677734375, output=1.3727264183
			11'd202: out = 32'b00000000000000001010111110010101; // input=0.19775390625, output=1.37173028174
			11'd203: out = 32'b00000000000000001010111101110100; // input=0.19873046875, output=1.37073394497
			11'd204: out = 32'b00000000000000001010111101010100; // input=0.19970703125, output=1.36973740686
			11'd205: out = 32'b00000000000000001010111100110011; // input=0.20068359375, output=1.36874066631
			11'd206: out = 32'b00000000000000001010111100010010; // input=0.20166015625, output=1.3677437222
			11'd207: out = 32'b00000000000000001010111011110010; // input=0.20263671875, output=1.36674657341
			11'd208: out = 32'b00000000000000001010111011010001; // input=0.20361328125, output=1.36574921883
			11'd209: out = 32'b00000000000000001010111010110000; // input=0.20458984375, output=1.36475165733
			11'd210: out = 32'b00000000000000001010111010001111; // input=0.20556640625, output=1.3637538878
			11'd211: out = 32'b00000000000000001010111001101111; // input=0.20654296875, output=1.36275590911
			11'd212: out = 32'b00000000000000001010111001001110; // input=0.20751953125, output=1.36175772013
			11'd213: out = 32'b00000000000000001010111000101101; // input=0.20849609375, output=1.36075931974
			11'd214: out = 32'b00000000000000001010111000001101; // input=0.20947265625, output=1.3597607068
			11'd215: out = 32'b00000000000000001010110111101100; // input=0.21044921875, output=1.35876188018
			11'd216: out = 32'b00000000000000001010110111001011; // input=0.21142578125, output=1.35776283875
			11'd217: out = 32'b00000000000000001010110110101010; // input=0.21240234375, output=1.35676358138
			11'd218: out = 32'b00000000000000001010110110001010; // input=0.21337890625, output=1.35576410692
			11'd219: out = 32'b00000000000000001010110101101001; // input=0.21435546875, output=1.35476441423
			11'd220: out = 32'b00000000000000001010110101001000; // input=0.21533203125, output=1.35376450217
			11'd221: out = 32'b00000000000000001010110100100111; // input=0.21630859375, output=1.35276436959
			11'd222: out = 32'b00000000000000001010110100000111; // input=0.21728515625, output=1.35176401536
			11'd223: out = 32'b00000000000000001010110011100110; // input=0.21826171875, output=1.35076343831
			11'd224: out = 32'b00000000000000001010110011000101; // input=0.21923828125, output=1.3497626373
			11'd225: out = 32'b00000000000000001010110010100100; // input=0.22021484375, output=1.34876161118
			11'd226: out = 32'b00000000000000001010110010000011; // input=0.22119140625, output=1.34776035878
			11'd227: out = 32'b00000000000000001010110001100011; // input=0.22216796875, output=1.34675887895
			11'd228: out = 32'b00000000000000001010110001000010; // input=0.22314453125, output=1.34575717054
			11'd229: out = 32'b00000000000000001010110000100001; // input=0.22412109375, output=1.34475523237
			11'd230: out = 32'b00000000000000001010110000000000; // input=0.22509765625, output=1.34375306328
			11'd231: out = 32'b00000000000000001010101111011111; // input=0.22607421875, output=1.34275066211
			11'd232: out = 32'b00000000000000001010101110111110; // input=0.22705078125, output=1.34174802769
			11'd233: out = 32'b00000000000000001010101110011110; // input=0.22802734375, output=1.34074515885
			11'd234: out = 32'b00000000000000001010101101111101; // input=0.22900390625, output=1.3397420544
			11'd235: out = 32'b00000000000000001010101101011100; // input=0.22998046875, output=1.33873871318
			11'd236: out = 32'b00000000000000001010101100111011; // input=0.23095703125, output=1.33773513401
			11'd237: out = 32'b00000000000000001010101100011010; // input=0.23193359375, output=1.3367313157
			11'd238: out = 32'b00000000000000001010101011111001; // input=0.23291015625, output=1.33572725708
			11'd239: out = 32'b00000000000000001010101011011000; // input=0.23388671875, output=1.33472295695
			11'd240: out = 32'b00000000000000001010101010110111; // input=0.23486328125, output=1.33371841413
			11'd241: out = 32'b00000000000000001010101010010110; // input=0.23583984375, output=1.33271362743
			11'd242: out = 32'b00000000000000001010101001110101; // input=0.23681640625, output=1.33170859566
			11'd243: out = 32'b00000000000000001010101001010100; // input=0.23779296875, output=1.33070331761
			11'd244: out = 32'b00000000000000001010101000110100; // input=0.23876953125, output=1.3296977921
			11'd245: out = 32'b00000000000000001010101000010011; // input=0.23974609375, output=1.32869201792
			11'd246: out = 32'b00000000000000001010100111110010; // input=0.24072265625, output=1.32768599387
			11'd247: out = 32'b00000000000000001010100111010001; // input=0.24169921875, output=1.32667971875
			11'd248: out = 32'b00000000000000001010100110110000; // input=0.24267578125, output=1.32567319134
			11'd249: out = 32'b00000000000000001010100110001111; // input=0.24365234375, output=1.32466641044
			11'd250: out = 32'b00000000000000001010100101101110; // input=0.24462890625, output=1.32365937483
			11'd251: out = 32'b00000000000000001010100101001101; // input=0.24560546875, output=1.3226520833
			11'd252: out = 32'b00000000000000001010100100101100; // input=0.24658203125, output=1.32164453463
			11'd253: out = 32'b00000000000000001010100100001011; // input=0.24755859375, output=1.3206367276
			11'd254: out = 32'b00000000000000001010100011101010; // input=0.24853515625, output=1.31962866098
			11'd255: out = 32'b00000000000000001010100011001001; // input=0.24951171875, output=1.31862033355
			11'd256: out = 32'b00000000000000001010100010101000; // input=0.25048828125, output=1.31761174409
			11'd257: out = 32'b00000000000000001010100010000110; // input=0.25146484375, output=1.31660289135
			11'd258: out = 32'b00000000000000001010100001100101; // input=0.25244140625, output=1.31559377412
			11'd259: out = 32'b00000000000000001010100001000100; // input=0.25341796875, output=1.31458439114
			11'd260: out = 32'b00000000000000001010100000100011; // input=0.25439453125, output=1.31357474118
			11'd261: out = 32'b00000000000000001010100000000010; // input=0.25537109375, output=1.312564823
			11'd262: out = 32'b00000000000000001010011111100001; // input=0.25634765625, output=1.31155463536
			11'd263: out = 32'b00000000000000001010011111000000; // input=0.25732421875, output=1.310544177
			11'd264: out = 32'b00000000000000001010011110011111; // input=0.25830078125, output=1.30953344668
			11'd265: out = 32'b00000000000000001010011101111110; // input=0.25927734375, output=1.30852244314
			11'd266: out = 32'b00000000000000001010011101011101; // input=0.26025390625, output=1.30751116513
			11'd267: out = 32'b00000000000000001010011100111011; // input=0.26123046875, output=1.30649961139
			11'd268: out = 32'b00000000000000001010011100011010; // input=0.26220703125, output=1.30548778065
			11'd269: out = 32'b00000000000000001010011011111001; // input=0.26318359375, output=1.30447567165
			11'd270: out = 32'b00000000000000001010011011011000; // input=0.26416015625, output=1.30346328313
			11'd271: out = 32'b00000000000000001010011010110111; // input=0.26513671875, output=1.30245061382
			11'd272: out = 32'b00000000000000001010011010010110; // input=0.26611328125, output=1.30143766244
			11'd273: out = 32'b00000000000000001010011001110100; // input=0.26708984375, output=1.30042442771
			11'd274: out = 32'b00000000000000001010011001010011; // input=0.26806640625, output=1.29941090836
			11'd275: out = 32'b00000000000000001010011000110010; // input=0.26904296875, output=1.2983971031
			11'd276: out = 32'b00000000000000001010011000010001; // input=0.27001953125, output=1.29738301066
			11'd277: out = 32'b00000000000000001010010111101111; // input=0.27099609375, output=1.29636862973
			11'd278: out = 32'b00000000000000001010010111001110; // input=0.27197265625, output=1.29535395904
			11'd279: out = 32'b00000000000000001010010110101101; // input=0.27294921875, output=1.29433899728
			11'd280: out = 32'b00000000000000001010010110001100; // input=0.27392578125, output=1.29332374316
			11'd281: out = 32'b00000000000000001010010101101010; // input=0.27490234375, output=1.29230819538
			11'd282: out = 32'b00000000000000001010010101001001; // input=0.27587890625, output=1.29129235264
			11'd283: out = 32'b00000000000000001010010100101000; // input=0.27685546875, output=1.29027621363
			11'd284: out = 32'b00000000000000001010010100000110; // input=0.27783203125, output=1.28925977704
			11'd285: out = 32'b00000000000000001010010011100101; // input=0.27880859375, output=1.28824304155
			11'd286: out = 32'b00000000000000001010010011000100; // input=0.27978515625, output=1.28722600586
			11'd287: out = 32'b00000000000000001010010010100010; // input=0.28076171875, output=1.28620866864
			11'd288: out = 32'b00000000000000001010010010000001; // input=0.28173828125, output=1.28519102857
			11'd289: out = 32'b00000000000000001010010001100000; // input=0.28271484375, output=1.28417308432
			11'd290: out = 32'b00000000000000001010010000111110; // input=0.28369140625, output=1.28315483458
			11'd291: out = 32'b00000000000000001010010000011101; // input=0.28466796875, output=1.28213627799
			11'd292: out = 32'b00000000000000001010001111111100; // input=0.28564453125, output=1.28111741324
			11'd293: out = 32'b00000000000000001010001111011010; // input=0.28662109375, output=1.28009823898
			11'd294: out = 32'b00000000000000001010001110111001; // input=0.28759765625, output=1.27907875386
			11'd295: out = 32'b00000000000000001010001110010111; // input=0.28857421875, output=1.27805895655
			11'd296: out = 32'b00000000000000001010001101110110; // input=0.28955078125, output=1.2770388457
			11'd297: out = 32'b00000000000000001010001101010101; // input=0.29052734375, output=1.27601841995
			11'd298: out = 32'b00000000000000001010001100110011; // input=0.29150390625, output=1.27499767795
			11'd299: out = 32'b00000000000000001010001100010010; // input=0.29248046875, output=1.27397661833
			11'd300: out = 32'b00000000000000001010001011110000; // input=0.29345703125, output=1.27295523974
			11'd301: out = 32'b00000000000000001010001011001111; // input=0.29443359375, output=1.27193354082
			11'd302: out = 32'b00000000000000001010001010101101; // input=0.29541015625, output=1.27091152019
			11'd303: out = 32'b00000000000000001010001010001100; // input=0.29638671875, output=1.26988917647
			11'd304: out = 32'b00000000000000001010001001101010; // input=0.29736328125, output=1.2688665083
			11'd305: out = 32'b00000000000000001010001001001001; // input=0.29833984375, output=1.2678435143
			11'd306: out = 32'b00000000000000001010001000100111; // input=0.29931640625, output=1.26682019307
			11'd307: out = 32'b00000000000000001010001000000110; // input=0.30029296875, output=1.26579654324
			11'd308: out = 32'b00000000000000001010000111100100; // input=0.30126953125, output=1.26477256342
			11'd309: out = 32'b00000000000000001010000111000011; // input=0.30224609375, output=1.2637482522
			11'd310: out = 32'b00000000000000001010000110100001; // input=0.30322265625, output=1.26272360819
			11'd311: out = 32'b00000000000000001010000101111111; // input=0.30419921875, output=1.26169863
			11'd312: out = 32'b00000000000000001010000101011110; // input=0.30517578125, output=1.2606733162
			11'd313: out = 32'b00000000000000001010000100111100; // input=0.30615234375, output=1.25964766541
			11'd314: out = 32'b00000000000000001010000100011011; // input=0.30712890625, output=1.2586216762
			11'd315: out = 32'b00000000000000001010000011111001; // input=0.30810546875, output=1.25759534715
			11'd316: out = 32'b00000000000000001010000011010111; // input=0.30908203125, output=1.25656867686
			11'd317: out = 32'b00000000000000001010000010110110; // input=0.31005859375, output=1.25554166389
			11'd318: out = 32'b00000000000000001010000010010100; // input=0.31103515625, output=1.25451430681
			11'd319: out = 32'b00000000000000001010000001110010; // input=0.31201171875, output=1.2534866042
			11'd320: out = 32'b00000000000000001010000001010001; // input=0.31298828125, output=1.25245855461
			11'd321: out = 32'b00000000000000001010000000101111; // input=0.31396484375, output=1.25143015662
			11'd322: out = 32'b00000000000000001010000000001101; // input=0.31494140625, output=1.25040140877
			11'd323: out = 32'b00000000000000001001111111101011; // input=0.31591796875, output=1.24937230962
			11'd324: out = 32'b00000000000000001001111111001010; // input=0.31689453125, output=1.24834285773
			11'd325: out = 32'b00000000000000001001111110101000; // input=0.31787109375, output=1.24731305162
			11'd326: out = 32'b00000000000000001001111110000110; // input=0.31884765625, output=1.24628288985
			11'd327: out = 32'b00000000000000001001111101100100; // input=0.31982421875, output=1.24525237094
			11'd328: out = 32'b00000000000000001001111101000011; // input=0.32080078125, output=1.24422149344
			11'd329: out = 32'b00000000000000001001111100100001; // input=0.32177734375, output=1.24319025588
			11'd330: out = 32'b00000000000000001001111011111111; // input=0.32275390625, output=1.24215865677
			11'd331: out = 32'b00000000000000001001111011011101; // input=0.32373046875, output=1.24112669464
			11'd332: out = 32'b00000000000000001001111010111011; // input=0.32470703125, output=1.240094368
			11'd333: out = 32'b00000000000000001001111010011010; // input=0.32568359375, output=1.23906167537
			11'd334: out = 32'b00000000000000001001111001111000; // input=0.32666015625, output=1.23802861525
			11'd335: out = 32'b00000000000000001001111001010110; // input=0.32763671875, output=1.23699518615
			11'd336: out = 32'b00000000000000001001111000110100; // input=0.32861328125, output=1.23596138656
			11'd337: out = 32'b00000000000000001001111000010010; // input=0.32958984375, output=1.23492721499
			11'd338: out = 32'b00000000000000001001110111110000; // input=0.33056640625, output=1.23389266992
			11'd339: out = 32'b00000000000000001001110111001110; // input=0.33154296875, output=1.23285774984
			11'd340: out = 32'b00000000000000001001110110101100; // input=0.33251953125, output=1.23182245324
			11'd341: out = 32'b00000000000000001001110110001010; // input=0.33349609375, output=1.23078677858
			11'd342: out = 32'b00000000000000001001110101101000; // input=0.33447265625, output=1.22975072435
			11'd343: out = 32'b00000000000000001001110101000111; // input=0.33544921875, output=1.228714289
			11'd344: out = 32'b00000000000000001001110100100101; // input=0.33642578125, output=1.22767747102
			11'd345: out = 32'b00000000000000001001110100000011; // input=0.33740234375, output=1.22664026885
			11'd346: out = 32'b00000000000000001001110011100001; // input=0.33837890625, output=1.22560268096
			11'd347: out = 32'b00000000000000001001110010111111; // input=0.33935546875, output=1.22456470579
			11'd348: out = 32'b00000000000000001001110010011101; // input=0.34033203125, output=1.22352634178
			11'd349: out = 32'b00000000000000001001110001111010; // input=0.34130859375, output=1.22248758739
			11'd350: out = 32'b00000000000000001001110001011000; // input=0.34228515625, output=1.22144844105
			11'd351: out = 32'b00000000000000001001110000110110; // input=0.34326171875, output=1.22040890119
			11'd352: out = 32'b00000000000000001001110000010100; // input=0.34423828125, output=1.21936896624
			11'd353: out = 32'b00000000000000001001101111110010; // input=0.34521484375, output=1.21832863463
			11'd354: out = 32'b00000000000000001001101111010000; // input=0.34619140625, output=1.21728790476
			11'd355: out = 32'b00000000000000001001101110101110; // input=0.34716796875, output=1.21624677506
			11'd356: out = 32'b00000000000000001001101110001100; // input=0.34814453125, output=1.21520524394
			11'd357: out = 32'b00000000000000001001101101101010; // input=0.34912109375, output=1.21416330979
			11'd358: out = 32'b00000000000000001001101101001000; // input=0.35009765625, output=1.21312097102
			11'd359: out = 32'b00000000000000001001101100100101; // input=0.35107421875, output=1.21207822602
			11'd360: out = 32'b00000000000000001001101100000011; // input=0.35205078125, output=1.21103507318
			11'd361: out = 32'b00000000000000001001101011100001; // input=0.35302734375, output=1.20999151089
			11'd362: out = 32'b00000000000000001001101010111111; // input=0.35400390625, output=1.20894753753
			11'd363: out = 32'b00000000000000001001101010011101; // input=0.35498046875, output=1.20790315147
			11'd364: out = 32'b00000000000000001001101001111010; // input=0.35595703125, output=1.20685835107
			11'd365: out = 32'b00000000000000001001101001011000; // input=0.35693359375, output=1.20581313471
			11'd366: out = 32'b00000000000000001001101000110110; // input=0.35791015625, output=1.20476750075
			11'd367: out = 32'b00000000000000001001101000010100; // input=0.35888671875, output=1.20372144753
			11'd368: out = 32'b00000000000000001001100111110001; // input=0.35986328125, output=1.20267497342
			11'd369: out = 32'b00000000000000001001100111001111; // input=0.36083984375, output=1.20162807674
			11'd370: out = 32'b00000000000000001001100110101101; // input=0.36181640625, output=1.20058075585
			11'd371: out = 32'b00000000000000001001100110001010; // input=0.36279296875, output=1.19953300907
			11'd372: out = 32'b00000000000000001001100101101000; // input=0.36376953125, output=1.19848483473
			11'd373: out = 32'b00000000000000001001100101000110; // input=0.36474609375, output=1.19743623116
			11'd374: out = 32'b00000000000000001001100100100011; // input=0.36572265625, output=1.19638719668
			11'd375: out = 32'b00000000000000001001100100000001; // input=0.36669921875, output=1.19533772959
			11'd376: out = 32'b00000000000000001001100011011110; // input=0.36767578125, output=1.19428782821
			11'd377: out = 32'b00000000000000001001100010111100; // input=0.36865234375, output=1.19323749083
			11'd378: out = 32'b00000000000000001001100010011010; // input=0.36962890625, output=1.19218671575
			11'd379: out = 32'b00000000000000001001100001110111; // input=0.37060546875, output=1.19113550126
			11'd380: out = 32'b00000000000000001001100001010101; // input=0.37158203125, output=1.19008384566
			11'd381: out = 32'b00000000000000001001100000110010; // input=0.37255859375, output=1.1890317472
			11'd382: out = 32'b00000000000000001001100000010000; // input=0.37353515625, output=1.18797920418
			11'd383: out = 32'b00000000000000001001011111101101; // input=0.37451171875, output=1.18692621486
			11'd384: out = 32'b00000000000000001001011111001011; // input=0.37548828125, output=1.18587277751
			11'd385: out = 32'b00000000000000001001011110101000; // input=0.37646484375, output=1.18481889037
			11'd386: out = 32'b00000000000000001001011110000110; // input=0.37744140625, output=1.1837645517
			11'd387: out = 32'b00000000000000001001011101100011; // input=0.37841796875, output=1.18270975975
			11'd388: out = 32'b00000000000000001001011101000000; // input=0.37939453125, output=1.18165451275
			11'd389: out = 32'b00000000000000001001011100011110; // input=0.38037109375, output=1.18059880895
			11'd390: out = 32'b00000000000000001001011011111011; // input=0.38134765625, output=1.17954264656
			11'd391: out = 32'b00000000000000001001011011011001; // input=0.38232421875, output=1.17848602382
			11'd392: out = 32'b00000000000000001001011010110110; // input=0.38330078125, output=1.17742893893
			11'd393: out = 32'b00000000000000001001011010010011; // input=0.38427734375, output=1.17637139011
			11'd394: out = 32'b00000000000000001001011001110001; // input=0.38525390625, output=1.17531337555
			11'd395: out = 32'b00000000000000001001011001001110; // input=0.38623046875, output=1.17425489347
			11'd396: out = 32'b00000000000000001001011000101011; // input=0.38720703125, output=1.17319594205
			11'd397: out = 32'b00000000000000001001011000001001; // input=0.38818359375, output=1.17213651948
			11'd398: out = 32'b00000000000000001001010111100110; // input=0.38916015625, output=1.17107662394
			11'd399: out = 32'b00000000000000001001010111000011; // input=0.39013671875, output=1.17001625359
			11'd400: out = 32'b00000000000000001001010110100000; // input=0.39111328125, output=1.16895540662
			11'd401: out = 32'b00000000000000001001010101111110; // input=0.39208984375, output=1.16789408118
			11'd402: out = 32'b00000000000000001001010101011011; // input=0.39306640625, output=1.16683227542
			11'd403: out = 32'b00000000000000001001010100111000; // input=0.39404296875, output=1.16576998749
			11'd404: out = 32'b00000000000000001001010100010101; // input=0.39501953125, output=1.16470721554
			11'd405: out = 32'b00000000000000001001010011110010; // input=0.39599609375, output=1.1636439577
			11'd406: out = 32'b00000000000000001001010011001111; // input=0.39697265625, output=1.16258021211
			11'd407: out = 32'b00000000000000001001010010101101; // input=0.39794921875, output=1.16151597687
			11'd408: out = 32'b00000000000000001001010010001010; // input=0.39892578125, output=1.16045125012
			11'd409: out = 32'b00000000000000001001010001100111; // input=0.39990234375, output=1.15938602995
			11'd410: out = 32'b00000000000000001001010001000100; // input=0.40087890625, output=1.15832031448
			11'd411: out = 32'b00000000000000001001010000100001; // input=0.40185546875, output=1.1572541018
			11'd412: out = 32'b00000000000000001001001111111110; // input=0.40283203125, output=1.15618738999
			11'd413: out = 32'b00000000000000001001001111011011; // input=0.40380859375, output=1.15512017715
			11'd414: out = 32'b00000000000000001001001110111000; // input=0.40478515625, output=1.15405246134
			11'd415: out = 32'b00000000000000001001001110010101; // input=0.40576171875, output=1.15298424064
			11'd416: out = 32'b00000000000000001001001101110010; // input=0.40673828125, output=1.15191551311
			11'd417: out = 32'b00000000000000001001001101001111; // input=0.40771484375, output=1.1508462768
			11'd418: out = 32'b00000000000000001001001100101100; // input=0.40869140625, output=1.14977652977
			11'd419: out = 32'b00000000000000001001001100001001; // input=0.40966796875, output=1.14870627005
			11'd420: out = 32'b00000000000000001001001011100110; // input=0.41064453125, output=1.14763549568
			11'd421: out = 32'b00000000000000001001001011000011; // input=0.41162109375, output=1.14656420469
			11'd422: out = 32'b00000000000000001001001010011111; // input=0.41259765625, output=1.14549239509
			11'd423: out = 32'b00000000000000001001001001111100; // input=0.41357421875, output=1.1444200649
			11'd424: out = 32'b00000000000000001001001001011001; // input=0.41455078125, output=1.14334721213
			11'd425: out = 32'b00000000000000001001001000110110; // input=0.41552734375, output=1.14227383477
			11'd426: out = 32'b00000000000000001001001000010011; // input=0.41650390625, output=1.14119993082
			11'd427: out = 32'b00000000000000001001000111110000; // input=0.41748046875, output=1.14012549826
			11'd428: out = 32'b00000000000000001001000111001100; // input=0.41845703125, output=1.13905053506
			11'd429: out = 32'b00000000000000001001000110101001; // input=0.41943359375, output=1.1379750392
			11'd430: out = 32'b00000000000000001001000110000110; // input=0.42041015625, output=1.13689900863
			11'd431: out = 32'b00000000000000001001000101100011; // input=0.42138671875, output=1.13582244131
			11'd432: out = 32'b00000000000000001001000100111111; // input=0.42236328125, output=1.13474533519
			11'd433: out = 32'b00000000000000001001000100011100; // input=0.42333984375, output=1.13366768821
			11'd434: out = 32'b00000000000000001001000011111001; // input=0.42431640625, output=1.13258949829
			11'd435: out = 32'b00000000000000001001000011010101; // input=0.42529296875, output=1.13151076336
			11'd436: out = 32'b00000000000000001001000010110010; // input=0.42626953125, output=1.13043148133
			11'd437: out = 32'b00000000000000001001000010001111; // input=0.42724609375, output=1.12935165012
			11'd438: out = 32'b00000000000000001001000001101011; // input=0.42822265625, output=1.12827126762
			11'd439: out = 32'b00000000000000001001000001001000; // input=0.42919921875, output=1.12719033172
			11'd440: out = 32'b00000000000000001001000000100100; // input=0.43017578125, output=1.12610884031
			11'd441: out = 32'b00000000000000001001000000000001; // input=0.43115234375, output=1.12502679127
			11'd442: out = 32'b00000000000000001000111111011101; // input=0.43212890625, output=1.12394418246
			11'd443: out = 32'b00000000000000001000111110111010; // input=0.43310546875, output=1.12286101173
			11'd444: out = 32'b00000000000000001000111110010110; // input=0.43408203125, output=1.12177727695
			11'd445: out = 32'b00000000000000001000111101110011; // input=0.43505859375, output=1.12069297596
			11'd446: out = 32'b00000000000000001000111101001111; // input=0.43603515625, output=1.11960810658
			11'd447: out = 32'b00000000000000001000111100101100; // input=0.43701171875, output=1.11852266665
			11'd448: out = 32'b00000000000000001000111100001000; // input=0.43798828125, output=1.11743665399
			11'd449: out = 32'b00000000000000001000111011100101; // input=0.43896484375, output=1.1163500664
			11'd450: out = 32'b00000000000000001000111011000001; // input=0.43994140625, output=1.11526290168
			11'd451: out = 32'b00000000000000001000111010011101; // input=0.44091796875, output=1.11417515763
			11'd452: out = 32'b00000000000000001000111001111010; // input=0.44189453125, output=1.11308683204
			11'd453: out = 32'b00000000000000001000111001010110; // input=0.44287109375, output=1.11199792267
			11'd454: out = 32'b00000000000000001000111000110010; // input=0.44384765625, output=1.11090842729
			11'd455: out = 32'b00000000000000001000111000001111; // input=0.44482421875, output=1.10981834366
			11'd456: out = 32'b00000000000000001000110111101011; // input=0.44580078125, output=1.10872766953
			11'd457: out = 32'b00000000000000001000110111000111; // input=0.44677734375, output=1.10763640264
			11'd458: out = 32'b00000000000000001000110110100011; // input=0.44775390625, output=1.10654454072
			11'd459: out = 32'b00000000000000001000110101111111; // input=0.44873046875, output=1.10545208149
			11'd460: out = 32'b00000000000000001000110101011100; // input=0.44970703125, output=1.10435902266
			11'd461: out = 32'b00000000000000001000110100111000; // input=0.45068359375, output=1.10326536194
			11'd462: out = 32'b00000000000000001000110100010100; // input=0.45166015625, output=1.10217109702
			11'd463: out = 32'b00000000000000001000110011110000; // input=0.45263671875, output=1.10107622559
			11'd464: out = 32'b00000000000000001000110011001100; // input=0.45361328125, output=1.09998074532
			11'd465: out = 32'b00000000000000001000110010101000; // input=0.45458984375, output=1.09888465389
			11'd466: out = 32'b00000000000000001000110010000100; // input=0.45556640625, output=1.09778794893
			11'd467: out = 32'b00000000000000001000110001100000; // input=0.45654296875, output=1.09669062811
			11'd468: out = 32'b00000000000000001000110000111100; // input=0.45751953125, output=1.09559268906
			11'd469: out = 32'b00000000000000001000110000011000; // input=0.45849609375, output=1.09449412941
			11'd470: out = 32'b00000000000000001000101111110100; // input=0.45947265625, output=1.09339494678
			11'd471: out = 32'b00000000000000001000101111010000; // input=0.46044921875, output=1.09229513877
			11'd472: out = 32'b00000000000000001000101110101100; // input=0.46142578125, output=1.09119470298
			11'd473: out = 32'b00000000000000001000101110001000; // input=0.46240234375, output=1.09009363702
			11'd474: out = 32'b00000000000000001000101101100100; // input=0.46337890625, output=1.08899193844
			11'd475: out = 32'b00000000000000001000101101000000; // input=0.46435546875, output=1.08788960482
			11'd476: out = 32'b00000000000000001000101100011100; // input=0.46533203125, output=1.08678663373
			11'd477: out = 32'b00000000000000001000101011111000; // input=0.46630859375, output=1.0856830227
			11'd478: out = 32'b00000000000000001000101011010011; // input=0.46728515625, output=1.08457876928
			11'd479: out = 32'b00000000000000001000101010101111; // input=0.46826171875, output=1.083473871
			11'd480: out = 32'b00000000000000001000101010001011; // input=0.46923828125, output=1.08236832536
			11'd481: out = 32'b00000000000000001000101001100111; // input=0.47021484375, output=1.08126212989
			11'd482: out = 32'b00000000000000001000101001000011; // input=0.47119140625, output=1.08015528208
			11'd483: out = 32'b00000000000000001000101000011110; // input=0.47216796875, output=1.07904777941
			11'd484: out = 32'b00000000000000001000100111111010; // input=0.47314453125, output=1.07793961935
			11'd485: out = 32'b00000000000000001000100111010110; // input=0.47412109375, output=1.07683079938
			11'd486: out = 32'b00000000000000001000100110110001; // input=0.47509765625, output=1.07572131695
			11'd487: out = 32'b00000000000000001000100110001101; // input=0.47607421875, output=1.0746111695
			11'd488: out = 32'b00000000000000001000100101101000; // input=0.47705078125, output=1.07350035446
			11'd489: out = 32'b00000000000000001000100101000100; // input=0.47802734375, output=1.07238886925
			11'd490: out = 32'b00000000000000001000100100100000; // input=0.47900390625, output=1.07127671129
			11'd491: out = 32'b00000000000000001000100011111011; // input=0.47998046875, output=1.07016387796
			11'd492: out = 32'b00000000000000001000100011010111; // input=0.48095703125, output=1.06905036667
			11'd493: out = 32'b00000000000000001000100010110010; // input=0.48193359375, output=1.06793617478
			11'd494: out = 32'b00000000000000001000100010001110; // input=0.48291015625, output=1.06682129967
			11'd495: out = 32'b00000000000000001000100001101001; // input=0.48388671875, output=1.06570573867
			11'd496: out = 32'b00000000000000001000100001000100; // input=0.48486328125, output=1.06458948915
			11'd497: out = 32'b00000000000000001000100000100000; // input=0.48583984375, output=1.06347254841
			11'd498: out = 32'b00000000000000001000011111111011; // input=0.48681640625, output=1.0623549138
			11'd499: out = 32'b00000000000000001000011111010111; // input=0.48779296875, output=1.0612365826
			11'd500: out = 32'b00000000000000001000011110110010; // input=0.48876953125, output=1.06011755212
			11'd501: out = 32'b00000000000000001000011110001101; // input=0.48974609375, output=1.05899781963
			11'd502: out = 32'b00000000000000001000011101101001; // input=0.49072265625, output=1.05787738241
			11'd503: out = 32'b00000000000000001000011101000100; // input=0.49169921875, output=1.05675623772
			11'd504: out = 32'b00000000000000001000011100011111; // input=0.49267578125, output=1.05563438281
			11'd505: out = 32'b00000000000000001000011011111010; // input=0.49365234375, output=1.0545118149
			11'd506: out = 32'b00000000000000001000011011010101; // input=0.49462890625, output=1.05338853122
			11'd507: out = 32'b00000000000000001000011010110001; // input=0.49560546875, output=1.05226452897
			11'd508: out = 32'b00000000000000001000011010001100; // input=0.49658203125, output=1.05113980536
			11'd509: out = 32'b00000000000000001000011001100111; // input=0.49755859375, output=1.05001435757
			11'd510: out = 32'b00000000000000001000011001000010; // input=0.49853515625, output=1.04888818277
			11'd511: out = 32'b00000000000000001000011000011101; // input=0.49951171875, output=1.04776127811
			11'd512: out = 32'b00000000000000001000010111111000; // input=0.50048828125, output=1.04663364075
			11'd513: out = 32'b00000000000000001000010111010011; // input=0.50146484375, output=1.04550526781
			11'd514: out = 32'b00000000000000001000010110101110; // input=0.50244140625, output=1.04437615641
			11'd515: out = 32'b00000000000000001000010110001001; // input=0.50341796875, output=1.04324630367
			11'd516: out = 32'b00000000000000001000010101100100; // input=0.50439453125, output=1.04211570666
			11'd517: out = 32'b00000000000000001000010100111111; // input=0.50537109375, output=1.04098436248
			11'd518: out = 32'b00000000000000001000010100011010; // input=0.50634765625, output=1.03985226819
			11'd519: out = 32'b00000000000000001000010011110101; // input=0.50732421875, output=1.03871942083
			11'd520: out = 32'b00000000000000001000010011010000; // input=0.50830078125, output=1.03758581745
			11'd521: out = 32'b00000000000000001000010010101010; // input=0.50927734375, output=1.03645145508
			11'd522: out = 32'b00000000000000001000010010000101; // input=0.51025390625, output=1.03531633071
			11'd523: out = 32'b00000000000000001000010001100000; // input=0.51123046875, output=1.03418044136
			11'd524: out = 32'b00000000000000001000010000111011; // input=0.51220703125, output=1.033043784
			11'd525: out = 32'b00000000000000001000010000010110; // input=0.51318359375, output=1.03190635561
			11'd526: out = 32'b00000000000000001000001111110000; // input=0.51416015625, output=1.03076815313
			11'd527: out = 32'b00000000000000001000001111001011; // input=0.51513671875, output=1.0296291735
			11'd528: out = 32'b00000000000000001000001110100110; // input=0.51611328125, output=1.02848941365
			11'd529: out = 32'b00000000000000001000001110000000; // input=0.51708984375, output=1.0273488705
			11'd530: out = 32'b00000000000000001000001101011011; // input=0.51806640625, output=1.02620754093
			11'd531: out = 32'b00000000000000001000001100110101; // input=0.51904296875, output=1.02506542184
			11'd532: out = 32'b00000000000000001000001100010000; // input=0.52001953125, output=1.02392251008
			11'd533: out = 32'b00000000000000001000001011101010; // input=0.52099609375, output=1.0227788025
			11'd534: out = 32'b00000000000000001000001011000101; // input=0.52197265625, output=1.02163429595
			11'd535: out = 32'b00000000000000001000001010011111; // input=0.52294921875, output=1.02048898724
			11'd536: out = 32'b00000000000000001000001001111010; // input=0.52392578125, output=1.01934287318
			11'd537: out = 32'b00000000000000001000001001010100; // input=0.52490234375, output=1.01819595056
			11'd538: out = 32'b00000000000000001000001000101111; // input=0.52587890625, output=1.01704821615
			11'd539: out = 32'b00000000000000001000001000001001; // input=0.52685546875, output=1.01589966671
			11'd540: out = 32'b00000000000000001000000111100011; // input=0.52783203125, output=1.01475029899
			11'd541: out = 32'b00000000000000001000000110111110; // input=0.52880859375, output=1.01360010971
			11'd542: out = 32'b00000000000000001000000110011000; // input=0.52978515625, output=1.01244909558
			11'd543: out = 32'b00000000000000001000000101110010; // input=0.53076171875, output=1.0112972533
			11'd544: out = 32'b00000000000000001000000101001100; // input=0.53173828125, output=1.01014457955
			11'd545: out = 32'b00000000000000001000000100100111; // input=0.53271484375, output=1.00899107098
			11'd546: out = 32'b00000000000000001000000100000001; // input=0.53369140625, output=1.00783672425
			11'd547: out = 32'b00000000000000001000000011011011; // input=0.53466796875, output=1.00668153598
			11'd548: out = 32'b00000000000000001000000010110101; // input=0.53564453125, output=1.00552550278
			11'd549: out = 32'b00000000000000001000000010001111; // input=0.53662109375, output=1.00436862125
			11'd550: out = 32'b00000000000000001000000001101001; // input=0.53759765625, output=1.00321088797
			11'd551: out = 32'b00000000000000001000000001000011; // input=0.53857421875, output=1.00205229949
			11'd552: out = 32'b00000000000000001000000000011101; // input=0.53955078125, output=1.00089285236
			11'd553: out = 32'b00000000000000000111111111110111; // input=0.54052734375, output=0.999732543114
			11'd554: out = 32'b00000000000000000111111111010001; // input=0.54150390625, output=0.998571368249
			11'd555: out = 32'b00000000000000000111111110101011; // input=0.54248046875, output=0.99740932426
			11'd556: out = 32'b00000000000000000111111110000101; // input=0.54345703125, output=0.996246407619
			11'd557: out = 32'b00000000000000000111111101011111; // input=0.54443359375, output=0.995082614781
			11'd558: out = 32'b00000000000000000111111100111001; // input=0.54541015625, output=0.993917942183
			11'd559: out = 32'b00000000000000000111111100010011; // input=0.54638671875, output=0.992752386243
			11'd560: out = 32'b00000000000000000111111011101100; // input=0.54736328125, output=0.991585943361
			11'd561: out = 32'b00000000000000000111111011000110; // input=0.54833984375, output=0.990418609919
			11'd562: out = 32'b00000000000000000111111010100000; // input=0.54931640625, output=0.989250382279
			11'd563: out = 32'b00000000000000000111111001111001; // input=0.55029296875, output=0.988081256785
			11'd564: out = 32'b00000000000000000111111001010011; // input=0.55126953125, output=0.986911229762
			11'd565: out = 32'b00000000000000000111111000101101; // input=0.55224609375, output=0.985740297517
			11'd566: out = 32'b00000000000000000111111000000110; // input=0.55322265625, output=0.984568456334
			11'd567: out = 32'b00000000000000000111110111100000; // input=0.55419921875, output=0.983395702482
			11'd568: out = 32'b00000000000000000111110110111001; // input=0.55517578125, output=0.982222032208
			11'd569: out = 32'b00000000000000000111110110010011; // input=0.55615234375, output=0.98104744174
			11'd570: out = 32'b00000000000000000111110101101100; // input=0.55712890625, output=0.979871927286
			11'd571: out = 32'b00000000000000000111110101000110; // input=0.55810546875, output=0.978695485033
			11'd572: out = 32'b00000000000000000111110100011111; // input=0.55908203125, output=0.977518111149
			11'd573: out = 32'b00000000000000000111110011111001; // input=0.56005859375, output=0.976339801781
			11'd574: out = 32'b00000000000000000111110011010010; // input=0.56103515625, output=0.975160553056
			11'd575: out = 32'b00000000000000000111110010101011; // input=0.56201171875, output=0.973980361079
			11'd576: out = 32'b00000000000000000111110010000101; // input=0.56298828125, output=0.972799221937
			11'd577: out = 32'b00000000000000000111110001011110; // input=0.56396484375, output=0.971617131693
			11'd578: out = 32'b00000000000000000111110000110111; // input=0.56494140625, output=0.97043408639
			11'd579: out = 32'b00000000000000000111110000010000; // input=0.56591796875, output=0.96925008205
			11'd580: out = 32'b00000000000000000111101111101010; // input=0.56689453125, output=0.968065114672
			11'd581: out = 32'b00000000000000000111101111000011; // input=0.56787109375, output=0.966879180235
			11'd582: out = 32'b00000000000000000111101110011100; // input=0.56884765625, output=0.965692274695
			11'd583: out = 32'b00000000000000000111101101110101; // input=0.56982421875, output=0.964504393987
			11'd584: out = 32'b00000000000000000111101101001110; // input=0.57080078125, output=0.963315534023
			11'd585: out = 32'b00000000000000000111101100100111; // input=0.57177734375, output=0.962125690692
			11'd586: out = 32'b00000000000000000111101100000000; // input=0.57275390625, output=0.960934859862
			11'd587: out = 32'b00000000000000000111101011011001; // input=0.57373046875, output=0.959743037376
			11'd588: out = 32'b00000000000000000111101010110010; // input=0.57470703125, output=0.958550219057
			11'd589: out = 32'b00000000000000000111101010001011; // input=0.57568359375, output=0.957356400702
			11'd590: out = 32'b00000000000000000111101001100100; // input=0.57666015625, output=0.956161578087
			11'd591: out = 32'b00000000000000000111101000111100; // input=0.57763671875, output=0.954965746961
			11'd592: out = 32'b00000000000000000111101000010101; // input=0.57861328125, output=0.953768903054
			11'd593: out = 32'b00000000000000000111100111101110; // input=0.57958984375, output=0.952571042068
			11'd594: out = 32'b00000000000000000111100111000111; // input=0.58056640625, output=0.951372159683
			11'd595: out = 32'b00000000000000000111100110011111; // input=0.58154296875, output=0.950172251554
			11'd596: out = 32'b00000000000000000111100101111000; // input=0.58251953125, output=0.948971313313
			11'd597: out = 32'b00000000000000000111100101010001; // input=0.58349609375, output=0.947769340563
			11'd598: out = 32'b00000000000000000111100100101001; // input=0.58447265625, output=0.946566328888
			11'd599: out = 32'b00000000000000000111100100000010; // input=0.58544921875, output=0.945362273841
			11'd600: out = 32'b00000000000000000111100011011010; // input=0.58642578125, output=0.944157170955
			11'd601: out = 32'b00000000000000000111100010110011; // input=0.58740234375, output=0.942951015732
			11'd602: out = 32'b00000000000000000111100010001011; // input=0.58837890625, output=0.941743803654
			11'd603: out = 32'b00000000000000000111100001100011; // input=0.58935546875, output=0.940535530172
			11'd604: out = 32'b00000000000000000111100000111100; // input=0.59033203125, output=0.939326190713
			11'd605: out = 32'b00000000000000000111100000010100; // input=0.59130859375, output=0.938115780679
			11'd606: out = 32'b00000000000000000111011111101100; // input=0.59228515625, output=0.936904295441
			11'd607: out = 32'b00000000000000000111011111000101; // input=0.59326171875, output=0.935691730348
			11'd608: out = 32'b00000000000000000111011110011101; // input=0.59423828125, output=0.934478080718
			11'd609: out = 32'b00000000000000000111011101110101; // input=0.59521484375, output=0.933263341845
			11'd610: out = 32'b00000000000000000111011101001101; // input=0.59619140625, output=0.932047508992
			11'd611: out = 32'b00000000000000000111011100100101; // input=0.59716796875, output=0.930830577396
			11'd612: out = 32'b00000000000000000111011011111110; // input=0.59814453125, output=0.929612542267
			11'd613: out = 32'b00000000000000000111011011010110; // input=0.59912109375, output=0.928393398785
			11'd614: out = 32'b00000000000000000111011010101110; // input=0.60009765625, output=0.9271731421
			11'd615: out = 32'b00000000000000000111011010000110; // input=0.60107421875, output=0.925951767338
			11'd616: out = 32'b00000000000000000111011001011110; // input=0.60205078125, output=0.924729269591
			11'd617: out = 32'b00000000000000000111011000110101; // input=0.60302734375, output=0.923505643923
			11'd618: out = 32'b00000000000000000111011000001101; // input=0.60400390625, output=0.922280885371
			11'd619: out = 32'b00000000000000000111010111100101; // input=0.60498046875, output=0.92105498894
			11'd620: out = 32'b00000000000000000111010110111101; // input=0.60595703125, output=0.919827949604
			11'd621: out = 32'b00000000000000000111010110010101; // input=0.60693359375, output=0.918599762308
			11'd622: out = 32'b00000000000000000111010101101100; // input=0.60791015625, output=0.917370421967
			11'd623: out = 32'b00000000000000000111010101000100; // input=0.60888671875, output=0.916139923464
			11'd624: out = 32'b00000000000000000111010100011100; // input=0.60986328125, output=0.91490826165
			11'd625: out = 32'b00000000000000000111010011110011; // input=0.61083984375, output=0.913675431347
			11'd626: out = 32'b00000000000000000111010011001011; // input=0.61181640625, output=0.912441427344
			11'd627: out = 32'b00000000000000000111010010100010; // input=0.61279296875, output=0.911206244396
			11'd628: out = 32'b00000000000000000111010001111010; // input=0.61376953125, output=0.90996987723
			11'd629: out = 32'b00000000000000000111010001010001; // input=0.61474609375, output=0.908732320536
			11'd630: out = 32'b00000000000000000111010000101001; // input=0.61572265625, output=0.907493568975
			11'd631: out = 32'b00000000000000000111010000000000; // input=0.61669921875, output=0.906253617171
			11'd632: out = 32'b00000000000000000111001111010111; // input=0.61767578125, output=0.905012459718
			11'd633: out = 32'b00000000000000000111001110101111; // input=0.61865234375, output=0.903770091174
			11'd634: out = 32'b00000000000000000111001110000110; // input=0.61962890625, output=0.902526506063
			11'd635: out = 32'b00000000000000000111001101011101; // input=0.62060546875, output=0.901281698877
			11'd636: out = 32'b00000000000000000111001100110100; // input=0.62158203125, output=0.90003566407
			11'd637: out = 32'b00000000000000000111001100001011; // input=0.62255859375, output=0.898788396062
			11'd638: out = 32'b00000000000000000111001011100011; // input=0.62353515625, output=0.89753988924
			11'd639: out = 32'b00000000000000000111001010111010; // input=0.62451171875, output=0.896290137952
			11'd640: out = 32'b00000000000000000111001010010001; // input=0.62548828125, output=0.895039136512
			11'd641: out = 32'b00000000000000000111001001101000; // input=0.62646484375, output=0.893786879197
			11'd642: out = 32'b00000000000000000111001000111111; // input=0.62744140625, output=0.892533360247
			11'd643: out = 32'b00000000000000000111001000010101; // input=0.62841796875, output=0.891278573866
			11'd644: out = 32'b00000000000000000111000111101100; // input=0.62939453125, output=0.89002251422
			11'd645: out = 32'b00000000000000000111000111000011; // input=0.63037109375, output=0.888765175437
			11'd646: out = 32'b00000000000000000111000110011010; // input=0.63134765625, output=0.887506551607
			11'd647: out = 32'b00000000000000000111000101110001; // input=0.63232421875, output=0.886246636783
			11'd648: out = 32'b00000000000000000111000101000111; // input=0.63330078125, output=0.884985424977
			11'd649: out = 32'b00000000000000000111000100011110; // input=0.63427734375, output=0.883722910163
			11'd650: out = 32'b00000000000000000111000011110100; // input=0.63525390625, output=0.882459086276
			11'd651: out = 32'b00000000000000000111000011001011; // input=0.63623046875, output=0.881193947211
			11'd652: out = 32'b00000000000000000111000010100001; // input=0.63720703125, output=0.879927486821
			11'd653: out = 32'b00000000000000000111000001111000; // input=0.63818359375, output=0.87865969892
			11'd654: out = 32'b00000000000000000111000001001110; // input=0.63916015625, output=0.877390577281
			11'd655: out = 32'b00000000000000000111000000100101; // input=0.64013671875, output=0.876120115634
			11'd656: out = 32'b00000000000000000110111111111011; // input=0.64111328125, output=0.87484830767
			11'd657: out = 32'b00000000000000000110111111010001; // input=0.64208984375, output=0.873575147036
			11'd658: out = 32'b00000000000000000110111110101000; // input=0.64306640625, output=0.872300627335
			11'd659: out = 32'b00000000000000000110111101111110; // input=0.64404296875, output=0.871024742129
			11'd660: out = 32'b00000000000000000110111101010100; // input=0.64501953125, output=0.869747484936
			11'd661: out = 32'b00000000000000000110111100101010; // input=0.64599609375, output=0.86846884923
			11'd662: out = 32'b00000000000000000110111100000000; // input=0.64697265625, output=0.867188828442
			11'd663: out = 32'b00000000000000000110111011010110; // input=0.64794921875, output=0.865907415954
			11'd664: out = 32'b00000000000000000110111010101100; // input=0.64892578125, output=0.864624605109
			11'd665: out = 32'b00000000000000000110111010000010; // input=0.64990234375, output=0.863340389199
			11'd666: out = 32'b00000000000000000110111001011000; // input=0.65087890625, output=0.862054761472
			11'd667: out = 32'b00000000000000000110111000101110; // input=0.65185546875, output=0.860767715131
			11'd668: out = 32'b00000000000000000110111000000011; // input=0.65283203125, output=0.859479243329
			11'd669: out = 32'b00000000000000000110110111011001; // input=0.65380859375, output=0.858189339174
			11'd670: out = 32'b00000000000000000110110110101111; // input=0.65478515625, output=0.856897995724
			11'd671: out = 32'b00000000000000000110110110000100; // input=0.65576171875, output=0.85560520599
			11'd672: out = 32'b00000000000000000110110101011010; // input=0.65673828125, output=0.854310962935
			11'd673: out = 32'b00000000000000000110110100110000; // input=0.65771484375, output=0.85301525947
			11'd674: out = 32'b00000000000000000110110100000101; // input=0.65869140625, output=0.851718088457
			11'd675: out = 32'b00000000000000000110110011011011; // input=0.65966796875, output=0.850419442709
			11'd676: out = 32'b00000000000000000110110010110000; // input=0.66064453125, output=0.849119314986
			11'd677: out = 32'b00000000000000000110110010000101; // input=0.66162109375, output=0.847817697999
			11'd678: out = 32'b00000000000000000110110001011011; // input=0.66259765625, output=0.846514584405
			11'd679: out = 32'b00000000000000000110110000110000; // input=0.66357421875, output=0.845209966809
			11'd680: out = 32'b00000000000000000110110000000101; // input=0.66455078125, output=0.843903837763
			11'd681: out = 32'b00000000000000000110101111011010; // input=0.66552734375, output=0.842596189766
			11'd682: out = 32'b00000000000000000110101110101111; // input=0.66650390625, output=0.841287015262
			11'd683: out = 32'b00000000000000000110101110000100; // input=0.66748046875, output=0.839976306642
			11'd684: out = 32'b00000000000000000110101101011001; // input=0.66845703125, output=0.838664056239
			11'd685: out = 32'b00000000000000000110101100101110; // input=0.66943359375, output=0.837350256332
			11'd686: out = 32'b00000000000000000110101100000011; // input=0.67041015625, output=0.836034899144
			11'd687: out = 32'b00000000000000000110101011011000; // input=0.67138671875, output=0.83471797684
			11'd688: out = 32'b00000000000000000110101010101101; // input=0.67236328125, output=0.833399481527
			11'd689: out = 32'b00000000000000000110101010000010; // input=0.67333984375, output=0.832079405255
			11'd690: out = 32'b00000000000000000110101001010110; // input=0.67431640625, output=0.830757740015
			11'd691: out = 32'b00000000000000000110101000101011; // input=0.67529296875, output=0.829434477737
			11'd692: out = 32'b00000000000000000110100111111111; // input=0.67626953125, output=0.828109610293
			11'd693: out = 32'b00000000000000000110100111010100; // input=0.67724609375, output=0.826783129494
			11'd694: out = 32'b00000000000000000110100110101001; // input=0.67822265625, output=0.825455027087
			11'd695: out = 32'b00000000000000000110100101111101; // input=0.67919921875, output=0.824125294761
			11'd696: out = 32'b00000000000000000110100101010001; // input=0.68017578125, output=0.82279392414
			11'd697: out = 32'b00000000000000000110100100100110; // input=0.68115234375, output=0.821460906784
			11'd698: out = 32'b00000000000000000110100011111010; // input=0.68212890625, output=0.820126234191
			11'd699: out = 32'b00000000000000000110100011001110; // input=0.68310546875, output=0.818789897792
			11'd700: out = 32'b00000000000000000110100010100010; // input=0.68408203125, output=0.817451888955
			11'd701: out = 32'b00000000000000000110100001110110; // input=0.68505859375, output=0.81611219898
			11'd702: out = 32'b00000000000000000110100001001010; // input=0.68603515625, output=0.814770819101
			11'd703: out = 32'b00000000000000000110100000011110; // input=0.68701171875, output=0.813427740483
			11'd704: out = 32'b00000000000000000110011111110010; // input=0.68798828125, output=0.812082954226
			11'd705: out = 32'b00000000000000000110011111000110; // input=0.68896484375, output=0.810736451356
			11'd706: out = 32'b00000000000000000110011110011010; // input=0.68994140625, output=0.809388222833
			11'd707: out = 32'b00000000000000000110011101101110; // input=0.69091796875, output=0.808038259545
			11'd708: out = 32'b00000000000000000110011101000010; // input=0.69189453125, output=0.806686552309
			11'd709: out = 32'b00000000000000000110011100010101; // input=0.69287109375, output=0.805333091869
			11'd710: out = 32'b00000000000000000110011011101001; // input=0.69384765625, output=0.803977868896
			11'd711: out = 32'b00000000000000000110011010111100; // input=0.69482421875, output=0.802620873988
			11'd712: out = 32'b00000000000000000110011010010000; // input=0.69580078125, output=0.801262097667
			11'd713: out = 32'b00000000000000000110011001100011; // input=0.69677734375, output=0.799901530381
			11'd714: out = 32'b00000000000000000110011000110111; // input=0.69775390625, output=0.798539162501
			11'd715: out = 32'b00000000000000000110011000001010; // input=0.69873046875, output=0.79717498432
			11'd716: out = 32'b00000000000000000110010111011101; // input=0.69970703125, output=0.795808986053
			11'd717: out = 32'b00000000000000000110010110110000; // input=0.70068359375, output=0.794441157837
			11'd718: out = 32'b00000000000000000110010110000011; // input=0.70166015625, output=0.793071489728
			11'd719: out = 32'b00000000000000000110010101010110; // input=0.70263671875, output=0.791699971702
			11'd720: out = 32'b00000000000000000110010100101001; // input=0.70361328125, output=0.790326593651
			11'd721: out = 32'b00000000000000000110010011111100; // input=0.70458984375, output=0.788951345388
			11'd722: out = 32'b00000000000000000110010011001111; // input=0.70556640625, output=0.787574216638
			11'd723: out = 32'b00000000000000000110010010100010; // input=0.70654296875, output=0.786195197045
			11'd724: out = 32'b00000000000000000110010001110101; // input=0.70751953125, output=0.784814276165
			11'd725: out = 32'b00000000000000000110010001000111; // input=0.70849609375, output=0.783431443467
			11'd726: out = 32'b00000000000000000110010000011010; // input=0.70947265625, output=0.782046688334
			11'd727: out = 32'b00000000000000000110001111101101; // input=0.71044921875, output=0.78066000006
			11'd728: out = 32'b00000000000000000110001110111111; // input=0.71142578125, output=0.779271367848
			11'd729: out = 32'b00000000000000000110001110010010; // input=0.71240234375, output=0.77788078081
			11'd730: out = 32'b00000000000000000110001101100100; // input=0.71337890625, output=0.776488227967
			11'd731: out = 32'b00000000000000000110001100110110; // input=0.71435546875, output=0.775093698247
			11'd732: out = 32'b00000000000000000110001100001001; // input=0.71533203125, output=0.773697180483
			11'd733: out = 32'b00000000000000000110001011011011; // input=0.71630859375, output=0.772298663413
			11'd734: out = 32'b00000000000000000110001010101101; // input=0.71728515625, output=0.770898135678
			11'd735: out = 32'b00000000000000000110001001111111; // input=0.71826171875, output=0.769495585822
			11'd736: out = 32'b00000000000000000110001001010001; // input=0.71923828125, output=0.768091002289
			11'd737: out = 32'b00000000000000000110001000100011; // input=0.72021484375, output=0.766684373425
			11'd738: out = 32'b00000000000000000110000111110101; // input=0.72119140625, output=0.765275687473
			11'd739: out = 32'b00000000000000000110000111000110; // input=0.72216796875, output=0.763864932573
			11'd740: out = 32'b00000000000000000110000110011000; // input=0.72314453125, output=0.762452096763
			11'd741: out = 32'b00000000000000000110000101101010; // input=0.72412109375, output=0.761037167974
			11'd742: out = 32'b00000000000000000110000100111011; // input=0.72509765625, output=0.759620134032
			11'd743: out = 32'b00000000000000000110000100001101; // input=0.72607421875, output=0.758200982654
			11'd744: out = 32'b00000000000000000110000011011110; // input=0.72705078125, output=0.756779701448
			11'd745: out = 32'b00000000000000000110000010110000; // input=0.72802734375, output=0.755356277913
			11'd746: out = 32'b00000000000000000110000010000001; // input=0.72900390625, output=0.753930699434
			11'd747: out = 32'b00000000000000000110000001010010; // input=0.72998046875, output=0.752502953285
			11'd748: out = 32'b00000000000000000110000000100011; // input=0.73095703125, output=0.751073026622
			11'd749: out = 32'b00000000000000000101111111110100; // input=0.73193359375, output=0.749640906488
			11'd750: out = 32'b00000000000000000101111111000101; // input=0.73291015625, output=0.748206579806
			11'd751: out = 32'b00000000000000000101111110010110; // input=0.73388671875, output=0.746770033382
			11'd752: out = 32'b00000000000000000101111101100111; // input=0.73486328125, output=0.745331253898
			11'd753: out = 32'b00000000000000000101111100111000; // input=0.73583984375, output=0.743890227917
			11'd754: out = 32'b00000000000000000101111100001001; // input=0.73681640625, output=0.742446941877
			11'd755: out = 32'b00000000000000000101111011011001; // input=0.73779296875, output=0.741001382088
			11'd756: out = 32'b00000000000000000101111010101010; // input=0.73876953125, output=0.739553534736
			11'd757: out = 32'b00000000000000000101111001111010; // input=0.73974609375, output=0.738103385877
			11'd758: out = 32'b00000000000000000101111001001011; // input=0.74072265625, output=0.736650921436
			11'd759: out = 32'b00000000000000000101111000011011; // input=0.74169921875, output=0.735196127207
			11'd760: out = 32'b00000000000000000101110111101011; // input=0.74267578125, output=0.733738988847
			11'd761: out = 32'b00000000000000000101110110111011; // input=0.74365234375, output=0.73227949188
			11'd762: out = 32'b00000000000000000101110110001011; // input=0.74462890625, output=0.730817621692
			11'd763: out = 32'b00000000000000000101110101011011; // input=0.74560546875, output=0.729353363528
			11'd764: out = 32'b00000000000000000101110100101011; // input=0.74658203125, output=0.727886702492
			11'd765: out = 32'b00000000000000000101110011111011; // input=0.74755859375, output=0.726417623546
			11'd766: out = 32'b00000000000000000101110011001011; // input=0.74853515625, output=0.724946111505
			11'd767: out = 32'b00000000000000000101110010011011; // input=0.74951171875, output=0.723472151039
			11'd768: out = 32'b00000000000000000101110001101010; // input=0.75048828125, output=0.721995726665
			11'd769: out = 32'b00000000000000000101110000111010; // input=0.75146484375, output=0.720516822751
			11'd770: out = 32'b00000000000000000101110000001001; // input=0.75244140625, output=0.719035423513
			11'd771: out = 32'b00000000000000000101101111011001; // input=0.75341796875, output=0.717551513008
			11'd772: out = 32'b00000000000000000101101110101000; // input=0.75439453125, output=0.716065075138
			11'd773: out = 32'b00000000000000000101101101110111; // input=0.75537109375, output=0.714576093643
			11'd774: out = 32'b00000000000000000101101101000110; // input=0.75634765625, output=0.713084552103
			11'd775: out = 32'b00000000000000000101101100010101; // input=0.75732421875, output=0.711590433931
			11'd776: out = 32'b00000000000000000101101011100100; // input=0.75830078125, output=0.710093722376
			11'd777: out = 32'b00000000000000000101101010110011; // input=0.75927734375, output=0.708594400515
			11'd778: out = 32'b00000000000000000101101010000010; // input=0.76025390625, output=0.707092451256
			11'd779: out = 32'b00000000000000000101101001010001; // input=0.76123046875, output=0.70558785733
			11'd780: out = 32'b00000000000000000101101000011111; // input=0.76220703125, output=0.704080601293
			11'd781: out = 32'b00000000000000000101100111101110; // input=0.76318359375, output=0.702570665524
			11'd782: out = 32'b00000000000000000101100110111100; // input=0.76416015625, output=0.701058032216
			11'd783: out = 32'b00000000000000000101100110001011; // input=0.76513671875, output=0.699542683381
			11'd784: out = 32'b00000000000000000101100101011001; // input=0.76611328125, output=0.698024600842
			11'd785: out = 32'b00000000000000000101100100100111; // input=0.76708984375, output=0.696503766233
			11'd786: out = 32'b00000000000000000101100011110101; // input=0.76806640625, output=0.694980160996
			11'd787: out = 32'b00000000000000000101100011000011; // input=0.76904296875, output=0.693453766377
			11'd788: out = 32'b00000000000000000101100010010001; // input=0.77001953125, output=0.691924563422
			11'd789: out = 32'b00000000000000000101100001011111; // input=0.77099609375, output=0.690392532978
			11'd790: out = 32'b00000000000000000101100000101100; // input=0.77197265625, output=0.688857655687
			11'd791: out = 32'b00000000000000000101011111111010; // input=0.77294921875, output=0.687319911983
			11'd792: out = 32'b00000000000000000101011111001000; // input=0.77392578125, output=0.685779282091
			11'd793: out = 32'b00000000000000000101011110010101; // input=0.77490234375, output=0.684235746018
			11'd794: out = 32'b00000000000000000101011101100010; // input=0.77587890625, output=0.68268928356
			11'd795: out = 32'b00000000000000000101011100110000; // input=0.77685546875, output=0.681139874289
			11'd796: out = 32'b00000000000000000101011011111101; // input=0.77783203125, output=0.679587497552
			11'd797: out = 32'b00000000000000000101011011001010; // input=0.77880859375, output=0.678032132473
			11'd798: out = 32'b00000000000000000101011010010111; // input=0.77978515625, output=0.676473757941
			11'd799: out = 32'b00000000000000000101011001100100; // input=0.78076171875, output=0.674912352614
			11'd800: out = 32'b00000000000000000101011000110000; // input=0.78173828125, output=0.67334789491
			11'd801: out = 32'b00000000000000000101010111111101; // input=0.78271484375, output=0.671780363006
			11'd802: out = 32'b00000000000000000101010111001001; // input=0.78369140625, output=0.670209734833
			11'd803: out = 32'b00000000000000000101010110010110; // input=0.78466796875, output=0.668635988073
			11'd804: out = 32'b00000000000000000101010101100010; // input=0.78564453125, output=0.667059100154
			11'd805: out = 32'b00000000000000000101010100101110; // input=0.78662109375, output=0.665479048247
			11'd806: out = 32'b00000000000000000101010011111011; // input=0.78759765625, output=0.663895809262
			11'd807: out = 32'b00000000000000000101010011000111; // input=0.78857421875, output=0.662309359842
			11'd808: out = 32'b00000000000000000101010010010010; // input=0.78955078125, output=0.660719676359
			11'd809: out = 32'b00000000000000000101010001011110; // input=0.79052734375, output=0.659126734912
			11'd810: out = 32'b00000000000000000101010000101010; // input=0.79150390625, output=0.657530511322
			11'd811: out = 32'b00000000000000000101001111110110; // input=0.79248046875, output=0.655930981122
			11'd812: out = 32'b00000000000000000101001111000001; // input=0.79345703125, output=0.654328119562
			11'd813: out = 32'b00000000000000000101001110001100; // input=0.79443359375, output=0.652721901594
			11'd814: out = 32'b00000000000000000101001101011000; // input=0.79541015625, output=0.651112301876
			11'd815: out = 32'b00000000000000000101001100100011; // input=0.79638671875, output=0.649499294759
			11'd816: out = 32'b00000000000000000101001011101110; // input=0.79736328125, output=0.647882854289
			11'd817: out = 32'b00000000000000000101001010111001; // input=0.79833984375, output=0.646262954198
			11'd818: out = 32'b00000000000000000101001010000100; // input=0.79931640625, output=0.644639567897
			11'd819: out = 32'b00000000000000000101001001001110; // input=0.80029296875, output=0.643012668475
			11'd820: out = 32'b00000000000000000101001000011001; // input=0.80126953125, output=0.64138222869
			11'd821: out = 32'b00000000000000000101000111100011; // input=0.80224609375, output=0.639748220967
			11'd822: out = 32'b00000000000000000101000110101110; // input=0.80322265625, output=0.638110617386
			11'd823: out = 32'b00000000000000000101000101111000; // input=0.80419921875, output=0.636469389683
			11'd824: out = 32'b00000000000000000101000101000010; // input=0.80517578125, output=0.634824509238
			11'd825: out = 32'b00000000000000000101000100001100; // input=0.80615234375, output=0.633175947074
			11'd826: out = 32'b00000000000000000101000011010110; // input=0.80712890625, output=0.631523673845
			11'd827: out = 32'b00000000000000000101000010100000; // input=0.80810546875, output=0.629867659836
			11'd828: out = 32'b00000000000000000101000001101001; // input=0.80908203125, output=0.62820787495
			11'd829: out = 32'b00000000000000000101000000110011; // input=0.81005859375, output=0.626544288707
			11'd830: out = 32'b00000000000000000100111111111100; // input=0.81103515625, output=0.62487687023
			11'd831: out = 32'b00000000000000000100111111000101; // input=0.81201171875, output=0.623205588247
			11'd832: out = 32'b00000000000000000100111110001110; // input=0.81298828125, output=0.621530411074
			11'd833: out = 32'b00000000000000000100111101010111; // input=0.81396484375, output=0.619851306615
			11'd834: out = 32'b00000000000000000100111100100000; // input=0.81494140625, output=0.61816824235
			11'd835: out = 32'b00000000000000000100111011101001; // input=0.81591796875, output=0.616481185331
			11'd836: out = 32'b00000000000000000100111010110001; // input=0.81689453125, output=0.614790102169
			11'd837: out = 32'b00000000000000000100111001111010; // input=0.81787109375, output=0.61309495903
			11'd838: out = 32'b00000000000000000100111001000010; // input=0.81884765625, output=0.611395721625
			11'd839: out = 32'b00000000000000000100111000001010; // input=0.81982421875, output=0.6096923552
			11'd840: out = 32'b00000000000000000100110111010010; // input=0.82080078125, output=0.607984824531
			11'd841: out = 32'b00000000000000000100110110011010; // input=0.82177734375, output=0.60627309391
			11'd842: out = 32'b00000000000000000100110101100010; // input=0.82275390625, output=0.60455712714
			11'd843: out = 32'b00000000000000000100110100101010; // input=0.82373046875, output=0.602836887524
			11'd844: out = 32'b00000000000000000100110011110001; // input=0.82470703125, output=0.601112337854
			11'd845: out = 32'b00000000000000000100110010111001; // input=0.82568359375, output=0.599383440402
			11'd846: out = 32'b00000000000000000100110010000000; // input=0.82666015625, output=0.597650156911
			11'd847: out = 32'b00000000000000000100110001000111; // input=0.82763671875, output=0.595912448581
			11'd848: out = 32'b00000000000000000100110000001110; // input=0.82861328125, output=0.594170276064
			11'd849: out = 32'b00000000000000000100101111010101; // input=0.82958984375, output=0.592423599447
			11'd850: out = 32'b00000000000000000100101110011011; // input=0.83056640625, output=0.590672378243
			11'd851: out = 32'b00000000000000000100101101100010; // input=0.83154296875, output=0.588916571382
			11'd852: out = 32'b00000000000000000100101100101000; // input=0.83251953125, output=0.587156137194
			11'd853: out = 32'b00000000000000000100101011101110; // input=0.83349609375, output=0.585391033401
			11'd854: out = 32'b00000000000000000100101010110100; // input=0.83447265625, output=0.583621217101
			11'd855: out = 32'b00000000000000000100101001111010; // input=0.83544921875, output=0.58184664476
			11'd856: out = 32'b00000000000000000100101001000000; // input=0.83642578125, output=0.580067272194
			11'd857: out = 32'b00000000000000000100101000000101; // input=0.83740234375, output=0.578283054556
			11'd858: out = 32'b00000000000000000100100111001011; // input=0.83837890625, output=0.576493946324
			11'd859: out = 32'b00000000000000000100100110010000; // input=0.83935546875, output=0.574699901288
			11'd860: out = 32'b00000000000000000100100101010101; // input=0.84033203125, output=0.572900872529
			11'd861: out = 32'b00000000000000000100100100011010; // input=0.84130859375, output=0.571096812411
			11'd862: out = 32'b00000000000000000100100011011110; // input=0.84228515625, output=0.569287672562
			11'd863: out = 32'b00000000000000000100100010100011; // input=0.84326171875, output=0.567473403856
			11'd864: out = 32'b00000000000000000100100001100111; // input=0.84423828125, output=0.565653956402
			11'd865: out = 32'b00000000000000000100100000101100; // input=0.84521484375, output=0.563829279521
			11'd866: out = 32'b00000000000000000100011111110000; // input=0.84619140625, output=0.561999321734
			11'd867: out = 32'b00000000000000000100011110110011; // input=0.84716796875, output=0.560164030741
			11'd868: out = 32'b00000000000000000100011101110111; // input=0.84814453125, output=0.558323353402
			11'd869: out = 32'b00000000000000000100011100111011; // input=0.84912109375, output=0.556477235721
			11'd870: out = 32'b00000000000000000100011011111110; // input=0.85009765625, output=0.554625622823
			11'd871: out = 32'b00000000000000000100011011000001; // input=0.85107421875, output=0.552768458938
			11'd872: out = 32'b00000000000000000100011010000100; // input=0.85205078125, output=0.550905687375
			11'd873: out = 32'b00000000000000000100011001000111; // input=0.85302734375, output=0.549037250506
			11'd874: out = 32'b00000000000000000100011000001001; // input=0.85400390625, output=0.547163089742
			11'd875: out = 32'b00000000000000000100010111001100; // input=0.85498046875, output=0.545283145509
			11'd876: out = 32'b00000000000000000100010110001110; // input=0.85595703125, output=0.543397357226
			11'd877: out = 32'b00000000000000000100010101010000; // input=0.85693359375, output=0.541505663281
			11'd878: out = 32'b00000000000000000100010100010010; // input=0.85791015625, output=0.539608001008
			11'd879: out = 32'b00000000000000000100010011010011; // input=0.85888671875, output=0.537704306657
			11'd880: out = 32'b00000000000000000100010010010101; // input=0.85986328125, output=0.535794515372
			11'd881: out = 32'b00000000000000000100010001010110; // input=0.86083984375, output=0.533878561162
			11'd882: out = 32'b00000000000000000100010000010111; // input=0.86181640625, output=0.531956376874
			11'd883: out = 32'b00000000000000000100001111011000; // input=0.86279296875, output=0.530027894162
			11'd884: out = 32'b00000000000000000100001110011001; // input=0.86376953125, output=0.528093043461
			11'd885: out = 32'b00000000000000000100001101011001; // input=0.86474609375, output=0.526151753951
			11'd886: out = 32'b00000000000000000100001100011001; // input=0.86572265625, output=0.524203953531
			11'd887: out = 32'b00000000000000000100001011011001; // input=0.86669921875, output=0.522249568781
			11'd888: out = 32'b00000000000000000100001010011001; // input=0.86767578125, output=0.520288524932
			11'd889: out = 32'b00000000000000000100001001011000; // input=0.86865234375, output=0.51832074583
			11'd890: out = 32'b00000000000000000100001000011000; // input=0.86962890625, output=0.516346153897
			11'd891: out = 32'b00000000000000000100000111010111; // input=0.87060546875, output=0.514364670098
			11'd892: out = 32'b00000000000000000100000110010110; // input=0.87158203125, output=0.5123762139
			11'd893: out = 32'b00000000000000000100000101010100; // input=0.87255859375, output=0.51038070323
			11'd894: out = 32'b00000000000000000100000100010011; // input=0.87353515625, output=0.508378054438
			11'd895: out = 32'b00000000000000000100000011010001; // input=0.87451171875, output=0.506368182252
			11'd896: out = 32'b00000000000000000100000010001111; // input=0.87548828125, output=0.504350999733
			11'd897: out = 32'b00000000000000000100000001001100; // input=0.87646484375, output=0.502326418228
			11'd898: out = 32'b00000000000000000100000000001010; // input=0.87744140625, output=0.500294347326
			11'd899: out = 32'b00000000000000000011111111000111; // input=0.87841796875, output=0.498254694808
			11'd900: out = 32'b00000000000000000011111110000100; // input=0.87939453125, output=0.496207366591
			11'd901: out = 32'b00000000000000000011111101000000; // input=0.88037109375, output=0.494152266683
			11'd902: out = 32'b00000000000000000011111011111101; // input=0.88134765625, output=0.492089297121
			11'd903: out = 32'b00000000000000000011111010111001; // input=0.88232421875, output=0.490018357918
			11'd904: out = 32'b00000000000000000011111001110101; // input=0.88330078125, output=0.487939347004
			11'd905: out = 32'b00000000000000000011111000110000; // input=0.88427734375, output=0.485852160163
			11'd906: out = 32'b00000000000000000011110111101100; // input=0.88525390625, output=0.483756690969
			11'd907: out = 32'b00000000000000000011110110100111; // input=0.88623046875, output=0.481652830723
			11'd908: out = 32'b00000000000000000011110101100010; // input=0.88720703125, output=0.479540468383
			11'd909: out = 32'b00000000000000000011110100011100; // input=0.88818359375, output=0.47741949049
			11'd910: out = 32'b00000000000000000011110011010110; // input=0.88916015625, output=0.475289781097
			11'd911: out = 32'b00000000000000000011110010010000; // input=0.89013671875, output=0.473151221691
			11'd912: out = 32'b00000000000000000011110001001010; // input=0.89111328125, output=0.471003691115
			11'd913: out = 32'b00000000000000000011110000000011; // input=0.89208984375, output=0.468847065479
			11'd914: out = 32'b00000000000000000011101110111100; // input=0.89306640625, output=0.46668121808
			11'd915: out = 32'b00000000000000000011101101110101; // input=0.89404296875, output=0.464506019307
			11'd916: out = 32'b00000000000000000011101100101101; // input=0.89501953125, output=0.462321336549
			11'd917: out = 32'b00000000000000000011101011100101; // input=0.89599609375, output=0.460127034094
			11'd918: out = 32'b00000000000000000011101010011101; // input=0.89697265625, output=0.457922973032
			11'd919: out = 32'b00000000000000000011101001010101; // input=0.89794921875, output=0.455709011145
			11'd920: out = 32'b00000000000000000011101000001100; // input=0.89892578125, output=0.453485002794
			11'd921: out = 32'b00000000000000000011100111000011; // input=0.89990234375, output=0.451250798807
			11'd922: out = 32'b00000000000000000011100101111001; // input=0.90087890625, output=0.449006246355
			11'd923: out = 32'b00000000000000000011100100101111; // input=0.90185546875, output=0.446751188828
			11'd924: out = 32'b00000000000000000011100011100101; // input=0.90283203125, output=0.444485465699
			11'd925: out = 32'b00000000000000000011100010011010; // input=0.90380859375, output=0.442208912389
			11'd926: out = 32'b00000000000000000011100001001111; // input=0.90478515625, output=0.439921360122
			11'd927: out = 32'b00000000000000000011100000000100; // input=0.90576171875, output=0.437622635771
			11'd928: out = 32'b00000000000000000011011110111000; // input=0.90673828125, output=0.435312561704
			11'd929: out = 32'b00000000000000000011011101101100; // input=0.90771484375, output=0.432990955614
			11'd930: out = 32'b00000000000000000011011100100000; // input=0.90869140625, output=0.430657630348
			11'd931: out = 32'b00000000000000000011011011010011; // input=0.90966796875, output=0.428312393723
			11'd932: out = 32'b00000000000000000011011010000110; // input=0.91064453125, output=0.425955048337
			11'd933: out = 32'b00000000000000000011011000111000; // input=0.91162109375, output=0.423585391365
			11'd934: out = 32'b00000000000000000011010111101010; // input=0.91259765625, output=0.421203214354
			11'd935: out = 32'b00000000000000000011010110011100; // input=0.91357421875, output=0.418808302995
			11'd936: out = 32'b00000000000000000011010101001101; // input=0.91455078125, output=0.416400436898
			11'd937: out = 32'b00000000000000000011010011111101; // input=0.91552734375, output=0.413979389341
			11'd938: out = 32'b00000000000000000011010010101110; // input=0.91650390625, output=0.411544927017
			11'd939: out = 32'b00000000000000000011010001011101; // input=0.91748046875, output=0.409096809761
			11'd940: out = 32'b00000000000000000011010000001101; // input=0.91845703125, output=0.406634790267
			11'd941: out = 32'b00000000000000000011001110111011; // input=0.91943359375, output=0.404158613784
			11'd942: out = 32'b00000000000000000011001101101010; // input=0.92041015625, output=0.401668017804
			11'd943: out = 32'b00000000000000000011001100011000; // input=0.92138671875, output=0.399162731721
			11'd944: out = 32'b00000000000000000011001011000101; // input=0.92236328125, output=0.396642476482
			11'd945: out = 32'b00000000000000000011001001110010; // input=0.92333984375, output=0.394106964214
			11'd946: out = 32'b00000000000000000011001000011111; // input=0.92431640625, output=0.391555897824
			11'd947: out = 32'b00000000000000000011000111001010; // input=0.92529296875, output=0.388988970587
			11'd948: out = 32'b00000000000000000011000101110110; // input=0.92626953125, output=0.386405865698
			11'd949: out = 32'b00000000000000000011000100100001; // input=0.92724609375, output=0.383806255807
			11'd950: out = 32'b00000000000000000011000011001011; // input=0.92822265625, output=0.381189802517
			11'd951: out = 32'b00000000000000000011000001110101; // input=0.92919921875, output=0.378556155859
			11'd952: out = 32'b00000000000000000011000000011110; // input=0.93017578125, output=0.375904953732
			11'd953: out = 32'b00000000000000000010111111000110; // input=0.93115234375, output=0.3732358213
			11'd954: out = 32'b00000000000000000010111101101110; // input=0.93212890625, output=0.370548370363
			11'd955: out = 32'b00000000000000000010111100010101; // input=0.93310546875, output=0.36784219868
			11'd956: out = 32'b00000000000000000010111010111100; // input=0.93408203125, output=0.365116889244
			11'd957: out = 32'b00000000000000000010111001100010; // input=0.93505859375, output=0.362372009518
			11'd958: out = 32'b00000000000000000010111000001000; // input=0.93603515625, output=0.359607110609
			11'd959: out = 32'b00000000000000000010110110101100; // input=0.93701171875, output=0.356821726393
			11'd960: out = 32'b00000000000000000010110101010000; // input=0.93798828125, output=0.354015372576
			11'd961: out = 32'b00000000000000000010110011110100; // input=0.93896484375, output=0.351187545683
			11'd962: out = 32'b00000000000000000010110010010110; // input=0.93994140625, output=0.348337721984
			11'd963: out = 32'b00000000000000000010110000111000; // input=0.94091796875, output=0.345465356329
			11'd964: out = 32'b00000000000000000010101111011001; // input=0.94189453125, output=0.34256988091
			11'd965: out = 32'b00000000000000000010101101111010; // input=0.94287109375, output=0.339650703915
			11'd966: out = 32'b00000000000000000010101100011001; // input=0.94384765625, output=0.336707208087
			11'd967: out = 32'b00000000000000000010101010111000; // input=0.94482421875, output=0.333738749167
			11'd968: out = 32'b00000000000000000010101001010110; // input=0.94580078125, output=0.330744654211
			11'd969: out = 32'b00000000000000000010100111110011; // input=0.94677734375, output=0.327724219773
			11'd970: out = 32'b00000000000000000010100110001111; // input=0.94775390625, output=0.324676709931
			11'd971: out = 32'b00000000000000000010100100101010; // input=0.94873046875, output=0.321601354156
			11'd972: out = 32'b00000000000000000010100011000101; // input=0.94970703125, output=0.318497344988
			11'd973: out = 32'b00000000000000000010100001011110; // input=0.95068359375, output=0.315363835514
			11'd974: out = 32'b00000000000000000010011111110110; // input=0.95166015625, output=0.312199936613
			11'd975: out = 32'b00000000000000000010011110001101; // input=0.95263671875, output=0.309004713959
			11'd976: out = 32'b00000000000000000010011100100100; // input=0.95361328125, output=0.305777184735
			11'd977: out = 32'b00000000000000000010011010111001; // input=0.95458984375, output=0.302516314039
			11'd978: out = 32'b00000000000000000010011001001101; // input=0.95556640625, output=0.299221010939
			11'd979: out = 32'b00000000000000000010010111100000; // input=0.95654296875, output=0.295890124136
			11'd980: out = 32'b00000000000000000010010101110001; // input=0.95751953125, output=0.292522437183
			11'd981: out = 32'b00000000000000000010010100000010; // input=0.95849609375, output=0.289116663208
			11'd982: out = 32'b00000000000000000010010010010001; // input=0.95947265625, output=0.285671439076
			11'd983: out = 32'b00000000000000000010010000011111; // input=0.96044921875, output=0.282185318912
			11'd984: out = 32'b00000000000000000010001110101011; // input=0.96142578125, output=0.278656766898
			11'd985: out = 32'b00000000000000000010001100110110; // input=0.96240234375, output=0.275084149249
			11'd986: out = 32'b00000000000000000010001010111111; // input=0.96337890625, output=0.271465725233
			11'd987: out = 32'b00000000000000000010001001000111; // input=0.96435546875, output=0.267799637122
			11'd988: out = 32'b00000000000000000010000111001110; // input=0.96533203125, output=0.264083898876
			11'd989: out = 32'b00000000000000000010000101010010; // input=0.96630859375, output=0.260316383399
			11'd990: out = 32'b00000000000000000010000011010101; // input=0.96728515625, output=0.256494808104
			11'd991: out = 32'b00000000000000000010000001010110; // input=0.96826171875, output=0.252616718532
			11'd992: out = 32'b00000000000000000001111111010101; // input=0.96923828125, output=0.248679469682
			11'd993: out = 32'b00000000000000000001111101010010; // input=0.97021484375, output=0.244680204644
			11'd994: out = 32'b00000000000000000001111011001100; // input=0.97119140625, output=0.240615830061
			11'd995: out = 32'b00000000000000000001111001000101; // input=0.97216796875, output=0.236482987801
			11'd996: out = 32'b00000000000000000001110110111011; // input=0.97314453125, output=0.232278022117
			11'd997: out = 32'b00000000000000000001110100101111; // input=0.97412109375, output=0.227996941384
			11'd998: out = 32'b00000000000000000001110010100000; // input=0.97509765625, output=0.223635373253
			11'd999: out = 32'b00000000000000000001110000001110; // input=0.97607421875, output=0.219188511821
			11'd1000: out = 32'b00000000000000000001101101111010; // input=0.97705078125, output=0.214651054972
			11'd1001: out = 32'b00000000000000000001101011100010; // input=0.97802734375, output=0.210017129581
			11'd1002: out = 32'b00000000000000000001101001000111; // input=0.97900390625, output=0.20528020156
			11'd1003: out = 32'b00000000000000000001100110101000; // input=0.97998046875, output=0.200432966839
			11'd1004: out = 32'b00000000000000000001100100000101; // input=0.98095703125, output=0.195467218063
			11'd1005: out = 32'b00000000000000000001100001011110; // input=0.98193359375, output=0.19037368008
			11'd1006: out = 32'b00000000000000000001011110110011; // input=0.98291015625, output=0.185141804779
			11'd1007: out = 32'b00000000000000000001011100000010; // input=0.98388671875, output=0.179759512289
			11'd1008: out = 32'b00000000000000000001011001001101; // input=0.98486328125, output=0.17421286033
			11'd1009: out = 32'b00000000000000000001010110010001; // input=0.98583984375, output=0.168485615729
			11'd1010: out = 32'b00000000000000000001010011001111; // input=0.98681640625, output=0.162558690208
			11'd1011: out = 32'b00000000000000000001010000000101; // input=0.98779296875, output=0.15640938387
			11'd1012: out = 32'b00000000000000000001001100110100; // input=0.98876953125, output=0.150010349655
			11'd1013: out = 32'b00000000000000000001001001011001; // input=0.98974609375, output=0.143328141623
			11'd1014: out = 32'b00000000000000000001000101110011; // input=0.99072265625, output=0.136321122325
			11'd1015: out = 32'b00000000000000000001000010000001; // input=0.99169921875, output=0.128936345273
			11'd1016: out = 32'b00000000000000000000111110000000; // input=0.99267578125, output=0.121104722866
			11'd1017: out = 32'b00000000000000000000111001101110; // input=0.99365234375, output=0.112733163685
			11'd1018: out = 32'b00000000000000000000110101000110; // input=0.99462890625, output=0.103690971223
			11'd1019: out = 32'b00000000000000000000110000000001; // input=0.99560546875, output=0.0937843662666
			11'd1020: out = 32'b00000000000000000000101010010110; // input=0.99658203125, output=0.0827032963273
			11'd1021: out = 32'b00000000000000000000100011110010; // input=0.99755859375, output=0.0698913486493
			11'd1022: out = 32'b00000000000000000000011011101110; // input=0.99853515625, output=0.0541331971646
			11'd1023: out = 32'b00000000000000000000010000000000; // input=0.99951171875, output=0.0312512717055
			11'd1024: out = 32'b00000000000000001100100100100000; // input=-0.00048828125, output=1.57128460806
			11'd1025: out = 32'b00000000000000001100100101000000; // input=-0.00146484375, output=1.57226117107
			11'd1026: out = 32'b00000000000000001100100101100000; // input=-0.00244140625, output=1.57323773547
			11'd1027: out = 32'b00000000000000001100100110000000; // input=-0.00341796875, output=1.5742143022
			11'd1028: out = 32'b00000000000000001100100110100000; // input=-0.00439453125, output=1.57519087219
			11'd1029: out = 32'b00000000000000001100100111000000; // input=-0.00537109375, output=1.57616744637
			11'd1030: out = 32'b00000000000000001100100111100000; // input=-0.00634765625, output=1.57714402567
			11'd1031: out = 32'b00000000000000001100101000000000; // input=-0.00732421875, output=1.57812061103
			11'd1032: out = 32'b00000000000000001100101000100000; // input=-0.00830078125, output=1.57909720337
			11'd1033: out = 32'b00000000000000001100101001000000; // input=-0.00927734375, output=1.58007380363
			11'd1034: out = 32'b00000000000000001100101001100000; // input=-0.01025390625, output=1.58105041274
			11'd1035: out = 32'b00000000000000001100101010000000; // input=-0.01123046875, output=1.58202703163
			11'd1036: out = 32'b00000000000000001100101010100000; // input=-0.01220703125, output=1.58300366123
			11'd1037: out = 32'b00000000000000001100101011000000; // input=-0.01318359375, output=1.58398030248
			11'd1038: out = 32'b00000000000000001100101011100000; // input=-0.01416015625, output=1.5849569563
			11'd1039: out = 32'b00000000000000001100101100000000; // input=-0.01513671875, output=1.58593362363
			11'd1040: out = 32'b00000000000000001100101100100000; // input=-0.01611328125, output=1.5869103054
			11'd1041: out = 32'b00000000000000001100101101000000; // input=-0.01708984375, output=1.58788700254
			11'd1042: out = 32'b00000000000000001100101101100000; // input=-0.01806640625, output=1.58886371599
			11'd1043: out = 32'b00000000000000001100101110000000; // input=-0.01904296875, output=1.58984044667
			11'd1044: out = 32'b00000000000000001100101110100000; // input=-0.02001953125, output=1.59081719553
			11'd1045: out = 32'b00000000000000001100101111000000; // input=-0.02099609375, output=1.59179396349
			11'd1046: out = 32'b00000000000000001100101111100000; // input=-0.02197265625, output=1.59277075149
			11'd1047: out = 32'b00000000000000001100110000000000; // input=-0.02294921875, output=1.59374756045
			11'd1048: out = 32'b00000000000000001100110000100000; // input=-0.02392578125, output=1.59472439132
			11'd1049: out = 32'b00000000000000001100110001000000; // input=-0.02490234375, output=1.59570124503
			11'd1050: out = 32'b00000000000000001100110001100000; // input=-0.02587890625, output=1.59667812251
			11'd1051: out = 32'b00000000000000001100110010000000; // input=-0.02685546875, output=1.59765502469
			11'd1052: out = 32'b00000000000000001100110010100000; // input=-0.02783203125, output=1.59863195252
			11'd1053: out = 32'b00000000000000001100110011000000; // input=-0.02880859375, output=1.59960890691
			11'd1054: out = 32'b00000000000000001100110011100000; // input=-0.02978515625, output=1.60058588882
			11'd1055: out = 32'b00000000000000001100110100000000; // input=-0.03076171875, output=1.60156289916
			11'd1056: out = 32'b00000000000000001100110100100000; // input=-0.03173828125, output=1.60253993889
			11'd1057: out = 32'b00000000000000001100110101000000; // input=-0.03271484375, output=1.60351700893
			11'd1058: out = 32'b00000000000000001100110101100000; // input=-0.03369140625, output=1.60449411022
			11'd1059: out = 32'b00000000000000001100110110000000; // input=-0.03466796875, output=1.60547124369
			11'd1060: out = 32'b00000000000000001100110110100000; // input=-0.03564453125, output=1.60644841029
			11'd1061: out = 32'b00000000000000001100110111000000; // input=-0.03662109375, output=1.60742561094
			11'd1062: out = 32'b00000000000000001100110111100000; // input=-0.03759765625, output=1.60840284659
			11'd1063: out = 32'b00000000000000001100111000000000; // input=-0.03857421875, output=1.60938011817
			11'd1064: out = 32'b00000000000000001100111000100000; // input=-0.03955078125, output=1.61035742662
			11'd1065: out = 32'b00000000000000001100111001000000; // input=-0.04052734375, output=1.61133477288
			11'd1066: out = 32'b00000000000000001100111001100000; // input=-0.04150390625, output=1.61231215788
			11'd1067: out = 32'b00000000000000001100111010000000; // input=-0.04248046875, output=1.61328958257
			11'd1068: out = 32'b00000000000000001100111010100000; // input=-0.04345703125, output=1.61426704788
			11'd1069: out = 32'b00000000000000001100111011000000; // input=-0.04443359375, output=1.61524455475
			11'd1070: out = 32'b00000000000000001100111011100000; // input=-0.04541015625, output=1.61622210412
			11'd1071: out = 32'b00000000000000001100111100000000; // input=-0.04638671875, output=1.61719969694
			11'd1072: out = 32'b00000000000000001100111100100000; // input=-0.04736328125, output=1.61817733413
			11'd1073: out = 32'b00000000000000001100111101000000; // input=-0.04833984375, output=1.61915501665
			11'd1074: out = 32'b00000000000000001100111101100001; // input=-0.04931640625, output=1.62013274543
			11'd1075: out = 32'b00000000000000001100111110000001; // input=-0.05029296875, output=1.62111052141
			11'd1076: out = 32'b00000000000000001100111110100001; // input=-0.05126953125, output=1.62208834554
			11'd1077: out = 32'b00000000000000001100111111000001; // input=-0.05224609375, output=1.62306621875
			11'd1078: out = 32'b00000000000000001100111111100001; // input=-0.05322265625, output=1.624044142
			11'd1079: out = 32'b00000000000000001101000000000001; // input=-0.05419921875, output=1.62502211622
			11'd1080: out = 32'b00000000000000001101000000100001; // input=-0.05517578125, output=1.62600014235
			11'd1081: out = 32'b00000000000000001101000001000001; // input=-0.05615234375, output=1.62697822135
			11'd1082: out = 32'b00000000000000001101000001100001; // input=-0.05712890625, output=1.62795635416
			11'd1083: out = 32'b00000000000000001101000010000001; // input=-0.05810546875, output=1.62893454171
			11'd1084: out = 32'b00000000000000001101000010100001; // input=-0.05908203125, output=1.62991278496
			11'd1085: out = 32'b00000000000000001101000011000001; // input=-0.06005859375, output=1.63089108485
			11'd1086: out = 32'b00000000000000001101000011100001; // input=-0.06103515625, output=1.63186944233
			11'd1087: out = 32'b00000000000000001101000100000001; // input=-0.06201171875, output=1.63284785834
			11'd1088: out = 32'b00000000000000001101000100100001; // input=-0.06298828125, output=1.63382633383
			11'd1089: out = 32'b00000000000000001101000101000001; // input=-0.06396484375, output=1.63480486976
			11'd1090: out = 32'b00000000000000001101000101100001; // input=-0.06494140625, output=1.63578346706
			11'd1091: out = 32'b00000000000000001101000110000001; // input=-0.06591796875, output=1.63676212669
			11'd1092: out = 32'b00000000000000001101000110100001; // input=-0.06689453125, output=1.63774084959
			11'd1093: out = 32'b00000000000000001101000111000010; // input=-0.06787109375, output=1.63871963672
			11'd1094: out = 32'b00000000000000001101000111100010; // input=-0.06884765625, output=1.63969848903
			11'd1095: out = 32'b00000000000000001101001000000010; // input=-0.06982421875, output=1.64067740747
			11'd1096: out = 32'b00000000000000001101001000100010; // input=-0.07080078125, output=1.64165639298
			11'd1097: out = 32'b00000000000000001101001001000010; // input=-0.07177734375, output=1.64263544653
			11'd1098: out = 32'b00000000000000001101001001100010; // input=-0.07275390625, output=1.64361456906
			11'd1099: out = 32'b00000000000000001101001010000010; // input=-0.07373046875, output=1.64459376153
			11'd1100: out = 32'b00000000000000001101001010100010; // input=-0.07470703125, output=1.6455730249
			11'd1101: out = 32'b00000000000000001101001011000010; // input=-0.07568359375, output=1.64655236011
			11'd1102: out = 32'b00000000000000001101001011100010; // input=-0.07666015625, output=1.64753176812
			11'd1103: out = 32'b00000000000000001101001100000010; // input=-0.07763671875, output=1.64851124989
			11'd1104: out = 32'b00000000000000001101001100100011; // input=-0.07861328125, output=1.64949080637
			11'd1105: out = 32'b00000000000000001101001101000011; // input=-0.07958984375, output=1.65047043853
			11'd1106: out = 32'b00000000000000001101001101100011; // input=-0.08056640625, output=1.65145014731
			11'd1107: out = 32'b00000000000000001101001110000011; // input=-0.08154296875, output=1.65242993369
			11'd1108: out = 32'b00000000000000001101001110100011; // input=-0.08251953125, output=1.65340979861
			11'd1109: out = 32'b00000000000000001101001111000011; // input=-0.08349609375, output=1.65438974304
			11'd1110: out = 32'b00000000000000001101001111100011; // input=-0.08447265625, output=1.65536976794
			11'd1111: out = 32'b00000000000000001101010000000011; // input=-0.08544921875, output=1.65634987426
			11'd1112: out = 32'b00000000000000001101010000100011; // input=-0.08642578125, output=1.65733006298
			11'd1113: out = 32'b00000000000000001101010001000100; // input=-0.08740234375, output=1.65831033506
			11'd1114: out = 32'b00000000000000001101010001100100; // input=-0.08837890625, output=1.65929069145
			11'd1115: out = 32'b00000000000000001101010010000100; // input=-0.08935546875, output=1.66027113312
			11'd1116: out = 32'b00000000000000001101010010100100; // input=-0.09033203125, output=1.66125166104
			11'd1117: out = 32'b00000000000000001101010011000100; // input=-0.09130859375, output=1.66223227617
			11'd1118: out = 32'b00000000000000001101010011100100; // input=-0.09228515625, output=1.66321297948
			11'd1119: out = 32'b00000000000000001101010100000100; // input=-0.09326171875, output=1.66419377194
			11'd1120: out = 32'b00000000000000001101010100100100; // input=-0.09423828125, output=1.66517465451
			11'd1121: out = 32'b00000000000000001101010101000101; // input=-0.09521484375, output=1.66615562817
			11'd1122: out = 32'b00000000000000001101010101100101; // input=-0.09619140625, output=1.66713669388
			11'd1123: out = 32'b00000000000000001101010110000101; // input=-0.09716796875, output=1.66811785261
			11'd1124: out = 32'b00000000000000001101010110100101; // input=-0.09814453125, output=1.66909910534
			11'd1125: out = 32'b00000000000000001101010111000101; // input=-0.09912109375, output=1.67008045303
			11'd1126: out = 32'b00000000000000001101010111100101; // input=-0.10009765625, output=1.67106189666
			11'd1127: out = 32'b00000000000000001101011000000110; // input=-0.10107421875, output=1.67204343721
			11'd1128: out = 32'b00000000000000001101011000100110; // input=-0.10205078125, output=1.67302507565
			11'd1129: out = 32'b00000000000000001101011001000110; // input=-0.10302734375, output=1.67400681295
			11'd1130: out = 32'b00000000000000001101011001100110; // input=-0.10400390625, output=1.67498865008
			11'd1131: out = 32'b00000000000000001101011010000110; // input=-0.10498046875, output=1.67597058804
			11'd1132: out = 32'b00000000000000001101011010100110; // input=-0.10595703125, output=1.67695262779
			11'd1133: out = 32'b00000000000000001101011011000111; // input=-0.10693359375, output=1.67793477032
			11'd1134: out = 32'b00000000000000001101011011100111; // input=-0.10791015625, output=1.6789170166
			11'd1135: out = 32'b00000000000000001101011100000111; // input=-0.10888671875, output=1.67989936762
			11'd1136: out = 32'b00000000000000001101011100100111; // input=-0.10986328125, output=1.68088182435
			11'd1137: out = 32'b00000000000000001101011101000111; // input=-0.11083984375, output=1.68186438778
			11'd1138: out = 32'b00000000000000001101011101101000; // input=-0.11181640625, output=1.6828470589
			11'd1139: out = 32'b00000000000000001101011110001000; // input=-0.11279296875, output=1.68382983868
			11'd1140: out = 32'b00000000000000001101011110101000; // input=-0.11376953125, output=1.68481272812
			11'd1141: out = 32'b00000000000000001101011111001000; // input=-0.11474609375, output=1.6857957282
			11'd1142: out = 32'b00000000000000001101011111101000; // input=-0.11572265625, output=1.6867788399
			11'd1143: out = 32'b00000000000000001101100000001001; // input=-0.11669921875, output=1.68776206423
			11'd1144: out = 32'b00000000000000001101100000101001; // input=-0.11767578125, output=1.68874540215
			11'd1145: out = 32'b00000000000000001101100001001001; // input=-0.11865234375, output=1.68972885468
			11'd1146: out = 32'b00000000000000001101100001101001; // input=-0.11962890625, output=1.69071242279
			11'd1147: out = 32'b00000000000000001101100010001001; // input=-0.12060546875, output=1.69169610749
			11'd1148: out = 32'b00000000000000001101100010101010; // input=-0.12158203125, output=1.69267990976
			11'd1149: out = 32'b00000000000000001101100011001010; // input=-0.12255859375, output=1.69366383059
			11'd1150: out = 32'b00000000000000001101100011101010; // input=-0.12353515625, output=1.69464787099
			11'd1151: out = 32'b00000000000000001101100100001010; // input=-0.12451171875, output=1.69563203196
			11'd1152: out = 32'b00000000000000001101100100101011; // input=-0.12548828125, output=1.69661631448
			11'd1153: out = 32'b00000000000000001101100101001011; // input=-0.12646484375, output=1.69760071956
			11'd1154: out = 32'b00000000000000001101100101101011; // input=-0.12744140625, output=1.6985852482
			11'd1155: out = 32'b00000000000000001101100110001100; // input=-0.12841796875, output=1.69956990141
			11'd1156: out = 32'b00000000000000001101100110101100; // input=-0.12939453125, output=1.70055468017
			11'd1157: out = 32'b00000000000000001101100111001100; // input=-0.13037109375, output=1.7015395855
			11'd1158: out = 32'b00000000000000001101100111101100; // input=-0.13134765625, output=1.70252461839
			11'd1159: out = 32'b00000000000000001101101000001101; // input=-0.13232421875, output=1.70350977987
			11'd1160: out = 32'b00000000000000001101101000101101; // input=-0.13330078125, output=1.70449507093
			11'd1161: out = 32'b00000000000000001101101001001101; // input=-0.13427734375, output=1.70548049257
			11'd1162: out = 32'b00000000000000001101101001101101; // input=-0.13525390625, output=1.70646604582
			11'd1163: out = 32'b00000000000000001101101010001110; // input=-0.13623046875, output=1.70745173168
			11'd1164: out = 32'b00000000000000001101101010101110; // input=-0.13720703125, output=1.70843755116
			11'd1165: out = 32'b00000000000000001101101011001110; // input=-0.13818359375, output=1.70942350528
			11'd1166: out = 32'b00000000000000001101101011101111; // input=-0.13916015625, output=1.71040959504
			11'd1167: out = 32'b00000000000000001101101100001111; // input=-0.14013671875, output=1.71139582147
			11'd1168: out = 32'b00000000000000001101101100101111; // input=-0.14111328125, output=1.71238218558
			11'd1169: out = 32'b00000000000000001101101101010000; // input=-0.14208984375, output=1.71336868839
			11'd1170: out = 32'b00000000000000001101101101110000; // input=-0.14306640625, output=1.71435533091
			11'd1171: out = 32'b00000000000000001101101110010000; // input=-0.14404296875, output=1.71534211417
			11'd1172: out = 32'b00000000000000001101101110110001; // input=-0.14501953125, output=1.7163290392
			11'd1173: out = 32'b00000000000000001101101111010001; // input=-0.14599609375, output=1.717316107
			11'd1174: out = 32'b00000000000000001101101111110001; // input=-0.14697265625, output=1.71830331861
			11'd1175: out = 32'b00000000000000001101110000010010; // input=-0.14794921875, output=1.71929067505
			11'd1176: out = 32'b00000000000000001101110000110010; // input=-0.14892578125, output=1.72027817735
			11'd1177: out = 32'b00000000000000001101110001010010; // input=-0.14990234375, output=1.72126582653
			11'd1178: out = 32'b00000000000000001101110001110011; // input=-0.15087890625, output=1.72225362364
			11'd1179: out = 32'b00000000000000001101110010010011; // input=-0.15185546875, output=1.72324156968
			11'd1180: out = 32'b00000000000000001101110010110100; // input=-0.15283203125, output=1.72422966571
			11'd1181: out = 32'b00000000000000001101110011010100; // input=-0.15380859375, output=1.72521791275
			11'd1182: out = 32'b00000000000000001101110011110100; // input=-0.15478515625, output=1.72620631183
			11'd1183: out = 32'b00000000000000001101110100010101; // input=-0.15576171875, output=1.727194864
			11'd1184: out = 32'b00000000000000001101110100110101; // input=-0.15673828125, output=1.72818357029
			11'd1185: out = 32'b00000000000000001101110101010110; // input=-0.15771484375, output=1.72917243174
			11'd1186: out = 32'b00000000000000001101110101110110; // input=-0.15869140625, output=1.73016144939
			11'd1187: out = 32'b00000000000000001101110110010110; // input=-0.15966796875, output=1.73115062428
			11'd1188: out = 32'b00000000000000001101110110110111; // input=-0.16064453125, output=1.73213995746
			11'd1189: out = 32'b00000000000000001101110111010111; // input=-0.16162109375, output=1.73312944996
			11'd1190: out = 32'b00000000000000001101110111111000; // input=-0.16259765625, output=1.73411910285
			11'd1191: out = 32'b00000000000000001101111000011000; // input=-0.16357421875, output=1.73510891715
			11'd1192: out = 32'b00000000000000001101111000111000; // input=-0.16455078125, output=1.73609889394
			11'd1193: out = 32'b00000000000000001101111001011001; // input=-0.16552734375, output=1.73708903424
			11'd1194: out = 32'b00000000000000001101111001111001; // input=-0.16650390625, output=1.73807933913
			11'd1195: out = 32'b00000000000000001101111010011010; // input=-0.16748046875, output=1.73906980964
			11'd1196: out = 32'b00000000000000001101111010111010; // input=-0.16845703125, output=1.74006044684
			11'd1197: out = 32'b00000000000000001101111011011011; // input=-0.16943359375, output=1.74105125178
			11'd1198: out = 32'b00000000000000001101111011111011; // input=-0.17041015625, output=1.74204222552
			11'd1199: out = 32'b00000000000000001101111100011100; // input=-0.17138671875, output=1.74303336913
			11'd1200: out = 32'b00000000000000001101111100111100; // input=-0.17236328125, output=1.74402468365
			11'd1201: out = 32'b00000000000000001101111101011101; // input=-0.17333984375, output=1.74501617017
			11'd1202: out = 32'b00000000000000001101111101111101; // input=-0.17431640625, output=1.74600782973
			11'd1203: out = 32'b00000000000000001101111110011110; // input=-0.17529296875, output=1.74699966341
			11'd1204: out = 32'b00000000000000001101111110111110; // input=-0.17626953125, output=1.74799167227
			11'd1205: out = 32'b00000000000000001101111111011111; // input=-0.17724609375, output=1.74898385739
			11'd1206: out = 32'b00000000000000001101111111111111; // input=-0.17822265625, output=1.74997621983
			11'd1207: out = 32'b00000000000000001110000000100000; // input=-0.17919921875, output=1.75096876068
			11'd1208: out = 32'b00000000000000001110000001000000; // input=-0.18017578125, output=1.75196148099
			11'd1209: out = 32'b00000000000000001110000001100001; // input=-0.18115234375, output=1.75295438186
			11'd1210: out = 32'b00000000000000001110000010000001; // input=-0.18212890625, output=1.75394746435
			11'd1211: out = 32'b00000000000000001110000010100010; // input=-0.18310546875, output=1.75494072955
			11'd1212: out = 32'b00000000000000001110000011000010; // input=-0.18408203125, output=1.75593417853
			11'd1213: out = 32'b00000000000000001110000011100011; // input=-0.18505859375, output=1.75692781239
			11'd1214: out = 32'b00000000000000001110000100000100; // input=-0.18603515625, output=1.7579216322
			11'd1215: out = 32'b00000000000000001110000100100100; // input=-0.18701171875, output=1.75891563906
			11'd1216: out = 32'b00000000000000001110000101000101; // input=-0.18798828125, output=1.75990983405
			11'd1217: out = 32'b00000000000000001110000101100101; // input=-0.18896484375, output=1.76090421826
			11'd1218: out = 32'b00000000000000001110000110000110; // input=-0.18994140625, output=1.76189879278
			11'd1219: out = 32'b00000000000000001110000110100110; // input=-0.19091796875, output=1.76289355871
			11'd1220: out = 32'b00000000000000001110000111000111; // input=-0.19189453125, output=1.76388851714
			11'd1221: out = 32'b00000000000000001110000111101000; // input=-0.19287109375, output=1.76488366917
			11'd1222: out = 32'b00000000000000001110001000001000; // input=-0.19384765625, output=1.7658790159
			11'd1223: out = 32'b00000000000000001110001000101001; // input=-0.19482421875, output=1.76687455842
			11'd1224: out = 32'b00000000000000001110001001001010; // input=-0.19580078125, output=1.76787029786
			11'd1225: out = 32'b00000000000000001110001001101010; // input=-0.19677734375, output=1.76886623529
			11'd1226: out = 32'b00000000000000001110001010001011; // input=-0.19775390625, output=1.76986237185
			11'd1227: out = 32'b00000000000000001110001010101011; // input=-0.19873046875, output=1.77085870862
			11'd1228: out = 32'b00000000000000001110001011001100; // input=-0.19970703125, output=1.77185524673
			11'd1229: out = 32'b00000000000000001110001011101101; // input=-0.20068359375, output=1.77285198728
			11'd1230: out = 32'b00000000000000001110001100001101; // input=-0.20166015625, output=1.77384893139
			11'd1231: out = 32'b00000000000000001110001100101110; // input=-0.20263671875, output=1.77484608018
			11'd1232: out = 32'b00000000000000001110001101001111; // input=-0.20361328125, output=1.77584343476
			11'd1233: out = 32'b00000000000000001110001101110000; // input=-0.20458984375, output=1.77684099626
			11'd1234: out = 32'b00000000000000001110001110010000; // input=-0.20556640625, output=1.77783876579
			11'd1235: out = 32'b00000000000000001110001110110001; // input=-0.20654296875, output=1.77883674448
			11'd1236: out = 32'b00000000000000001110001111010010; // input=-0.20751953125, output=1.77983493346
			11'd1237: out = 32'b00000000000000001110001111110010; // input=-0.20849609375, output=1.78083333385
			11'd1238: out = 32'b00000000000000001110010000010011; // input=-0.20947265625, output=1.78183194679
			11'd1239: out = 32'b00000000000000001110010000110100; // input=-0.21044921875, output=1.78283077341
			11'd1240: out = 32'b00000000000000001110010001010101; // input=-0.21142578125, output=1.78382981483
			11'd1241: out = 32'b00000000000000001110010001110101; // input=-0.21240234375, output=1.78482907221
			11'd1242: out = 32'b00000000000000001110010010010110; // input=-0.21337890625, output=1.78582854667
			11'd1243: out = 32'b00000000000000001110010010110111; // input=-0.21435546875, output=1.78682823936
			11'd1244: out = 32'b00000000000000001110010011011000; // input=-0.21533203125, output=1.78782815142
			11'd1245: out = 32'b00000000000000001110010011111000; // input=-0.21630859375, output=1.788828284
			11'd1246: out = 32'b00000000000000001110010100011001; // input=-0.21728515625, output=1.78982863823
			11'd1247: out = 32'b00000000000000001110010100111010; // input=-0.21826171875, output=1.79082921528
			11'd1248: out = 32'b00000000000000001110010101011011; // input=-0.21923828125, output=1.79183001629
			11'd1249: out = 32'b00000000000000001110010101111011; // input=-0.22021484375, output=1.79283104241
			11'd1250: out = 32'b00000000000000001110010110011100; // input=-0.22119140625, output=1.79383229481
			11'd1251: out = 32'b00000000000000001110010110111101; // input=-0.22216796875, output=1.79483377464
			11'd1252: out = 32'b00000000000000001110010111011110; // input=-0.22314453125, output=1.79583548305
			11'd1253: out = 32'b00000000000000001110010111111111; // input=-0.22412109375, output=1.79683742122
			11'd1254: out = 32'b00000000000000001110011000100000; // input=-0.22509765625, output=1.79783959031
			11'd1255: out = 32'b00000000000000001110011001000000; // input=-0.22607421875, output=1.79884199148
			11'd1256: out = 32'b00000000000000001110011001100001; // input=-0.22705078125, output=1.7998446259
			11'd1257: out = 32'b00000000000000001110011010000010; // input=-0.22802734375, output=1.80084749474
			11'd1258: out = 32'b00000000000000001110011010100011; // input=-0.22900390625, output=1.80185059919
			11'd1259: out = 32'b00000000000000001110011011000100; // input=-0.22998046875, output=1.80285394041
			11'd1260: out = 32'b00000000000000001110011011100101; // input=-0.23095703125, output=1.80385751958
			11'd1261: out = 32'b00000000000000001110011100000110; // input=-0.23193359375, output=1.80486133789
			11'd1262: out = 32'b00000000000000001110011100100111; // input=-0.23291015625, output=1.80586539651
			11'd1263: out = 32'b00000000000000001110011101001000; // input=-0.23388671875, output=1.80686969664
			11'd1264: out = 32'b00000000000000001110011101101000; // input=-0.23486328125, output=1.80787423946
			11'd1265: out = 32'b00000000000000001110011110001001; // input=-0.23583984375, output=1.80887902616
			11'd1266: out = 32'b00000000000000001110011110101010; // input=-0.23681640625, output=1.80988405793
			11'd1267: out = 32'b00000000000000001110011111001011; // input=-0.23779296875, output=1.81088933598
			11'd1268: out = 32'b00000000000000001110011111101100; // input=-0.23876953125, output=1.81189486149
			11'd1269: out = 32'b00000000000000001110100000001101; // input=-0.23974609375, output=1.81290063567
			11'd1270: out = 32'b00000000000000001110100000101110; // input=-0.24072265625, output=1.81390665972
			11'd1271: out = 32'b00000000000000001110100001001111; // input=-0.24169921875, output=1.81491293484
			11'd1272: out = 32'b00000000000000001110100001110000; // input=-0.24267578125, output=1.81591946225
			11'd1273: out = 32'b00000000000000001110100010010001; // input=-0.24365234375, output=1.81692624315
			11'd1274: out = 32'b00000000000000001110100010110010; // input=-0.24462890625, output=1.81793327876
			11'd1275: out = 32'b00000000000000001110100011010011; // input=-0.24560546875, output=1.81894057029
			11'd1276: out = 32'b00000000000000001110100011110100; // input=-0.24658203125, output=1.81994811896
			11'd1277: out = 32'b00000000000000001110100100010101; // input=-0.24755859375, output=1.82095592599
			11'd1278: out = 32'b00000000000000001110100100110110; // input=-0.24853515625, output=1.82196399261
			11'd1279: out = 32'b00000000000000001110100101010111; // input=-0.24951171875, output=1.82297232004
			11'd1280: out = 32'b00000000000000001110100101111000; // input=-0.25048828125, output=1.8239809095
			11'd1281: out = 32'b00000000000000001110100110011001; // input=-0.25146484375, output=1.82498976223
			11'd1282: out = 32'b00000000000000001110100110111010; // input=-0.25244140625, output=1.82599887947
			11'd1283: out = 32'b00000000000000001110100111011011; // input=-0.25341796875, output=1.82700826245
			11'd1284: out = 32'b00000000000000001110100111111100; // input=-0.25439453125, output=1.82801791241
			11'd1285: out = 32'b00000000000000001110101000011110; // input=-0.25537109375, output=1.82902783059
			11'd1286: out = 32'b00000000000000001110101000111111; // input=-0.25634765625, output=1.83003801823
			11'd1287: out = 32'b00000000000000001110101001100000; // input=-0.25732421875, output=1.83104847659
			11'd1288: out = 32'b00000000000000001110101010000001; // input=-0.25830078125, output=1.83205920691
			11'd1289: out = 32'b00000000000000001110101010100010; // input=-0.25927734375, output=1.83307021045
			11'd1290: out = 32'b00000000000000001110101011000011; // input=-0.26025390625, output=1.83408148846
			11'd1291: out = 32'b00000000000000001110101011100100; // input=-0.26123046875, output=1.8350930422
			11'd1292: out = 32'b00000000000000001110101100000101; // input=-0.26220703125, output=1.83610487294
			11'd1293: out = 32'b00000000000000001110101100100111; // input=-0.26318359375, output=1.83711698194
			11'd1294: out = 32'b00000000000000001110101101001000; // input=-0.26416015625, output=1.83812937046
			11'd1295: out = 32'b00000000000000001110101101101001; // input=-0.26513671875, output=1.83914203977
			11'd1296: out = 32'b00000000000000001110101110001010; // input=-0.26611328125, output=1.84015499115
			11'd1297: out = 32'b00000000000000001110101110101011; // input=-0.26708984375, output=1.84116822588
			11'd1298: out = 32'b00000000000000001110101111001101; // input=-0.26806640625, output=1.84218174523
			11'd1299: out = 32'b00000000000000001110101111101110; // input=-0.26904296875, output=1.84319555049
			11'd1300: out = 32'b00000000000000001110110000001111; // input=-0.27001953125, output=1.84420964293
			11'd1301: out = 32'b00000000000000001110110000110000; // input=-0.27099609375, output=1.84522402386
			11'd1302: out = 32'b00000000000000001110110001010010; // input=-0.27197265625, output=1.84623869455
			11'd1303: out = 32'b00000000000000001110110001110011; // input=-0.27294921875, output=1.84725365631
			11'd1304: out = 32'b00000000000000001110110010010100; // input=-0.27392578125, output=1.84826891043
			11'd1305: out = 32'b00000000000000001110110010110101; // input=-0.27490234375, output=1.84928445821
			11'd1306: out = 32'b00000000000000001110110011010111; // input=-0.27587890625, output=1.85030030095
			11'd1307: out = 32'b00000000000000001110110011111000; // input=-0.27685546875, output=1.85131643996
			11'd1308: out = 32'b00000000000000001110110100011001; // input=-0.27783203125, output=1.85233287655
			11'd1309: out = 32'b00000000000000001110110100111011; // input=-0.27880859375, output=1.85334961204
			11'd1310: out = 32'b00000000000000001110110101011100; // input=-0.27978515625, output=1.85436664773
			11'd1311: out = 32'b00000000000000001110110101111101; // input=-0.28076171875, output=1.85538398495
			11'd1312: out = 32'b00000000000000001110110110011111; // input=-0.28173828125, output=1.85640162502
			11'd1313: out = 32'b00000000000000001110110111000000; // input=-0.28271484375, output=1.85741956927
			11'd1314: out = 32'b00000000000000001110110111100001; // input=-0.28369140625, output=1.85843781901
			11'd1315: out = 32'b00000000000000001110111000000011; // input=-0.28466796875, output=1.8594563756
			11'd1316: out = 32'b00000000000000001110111000100100; // input=-0.28564453125, output=1.86047524035
			11'd1317: out = 32'b00000000000000001110111001000101; // input=-0.28662109375, output=1.86149441461
			11'd1318: out = 32'b00000000000000001110111001100111; // input=-0.28759765625, output=1.86251389973
			11'd1319: out = 32'b00000000000000001110111010001000; // input=-0.28857421875, output=1.86353369704
			11'd1320: out = 32'b00000000000000001110111010101010; // input=-0.28955078125, output=1.86455380789
			11'd1321: out = 32'b00000000000000001110111011001011; // input=-0.29052734375, output=1.86557423364
			11'd1322: out = 32'b00000000000000001110111011101101; // input=-0.29150390625, output=1.86659497564
			11'd1323: out = 32'b00000000000000001110111100001110; // input=-0.29248046875, output=1.86761603526
			11'd1324: out = 32'b00000000000000001110111100110000; // input=-0.29345703125, output=1.86863741384
			11'd1325: out = 32'b00000000000000001110111101010001; // input=-0.29443359375, output=1.86965911277
			11'd1326: out = 32'b00000000000000001110111101110010; // input=-0.29541015625, output=1.8706811334
			11'd1327: out = 32'b00000000000000001110111110010100; // input=-0.29638671875, output=1.87170347712
			11'd1328: out = 32'b00000000000000001110111110110101; // input=-0.29736328125, output=1.87272614528
			11'd1329: out = 32'b00000000000000001110111111010111; // input=-0.29833984375, output=1.87374913929
			11'd1330: out = 32'b00000000000000001110111111111001; // input=-0.29931640625, output=1.87477246052
			11'd1331: out = 32'b00000000000000001111000000011010; // input=-0.30029296875, output=1.87579611035
			11'd1332: out = 32'b00000000000000001111000000111100; // input=-0.30126953125, output=1.87682009017
			11'd1333: out = 32'b00000000000000001111000001011101; // input=-0.30224609375, output=1.87784440139
			11'd1334: out = 32'b00000000000000001111000001111111; // input=-0.30322265625, output=1.8788690454
			11'd1335: out = 32'b00000000000000001111000010100000; // input=-0.30419921875, output=1.87989402359
			11'd1336: out = 32'b00000000000000001111000011000010; // input=-0.30517578125, output=1.88091933739
			11'd1337: out = 32'b00000000000000001111000011100100; // input=-0.30615234375, output=1.88194498818
			11'd1338: out = 32'b00000000000000001111000100000101; // input=-0.30712890625, output=1.88297097739
			11'd1339: out = 32'b00000000000000001111000100100111; // input=-0.30810546875, output=1.88399730643
			11'd1340: out = 32'b00000000000000001111000101001000; // input=-0.30908203125, output=1.88502397673
			11'd1341: out = 32'b00000000000000001111000101101010; // input=-0.31005859375, output=1.8860509897
			11'd1342: out = 32'b00000000000000001111000110001100; // input=-0.31103515625, output=1.88707834678
			11'd1343: out = 32'b00000000000000001111000110101101; // input=-0.31201171875, output=1.88810604939
			11'd1344: out = 32'b00000000000000001111000111001111; // input=-0.31298828125, output=1.88913409898
			11'd1345: out = 32'b00000000000000001111000111110001; // input=-0.31396484375, output=1.89016249697
			11'd1346: out = 32'b00000000000000001111001000010011; // input=-0.31494140625, output=1.89119124482
			11'd1347: out = 32'b00000000000000001111001000110100; // input=-0.31591796875, output=1.89222034396
			11'd1348: out = 32'b00000000000000001111001001010110; // input=-0.31689453125, output=1.89324979586
			11'd1349: out = 32'b00000000000000001111001001111000; // input=-0.31787109375, output=1.89427960197
			11'd1350: out = 32'b00000000000000001111001010011010; // input=-0.31884765625, output=1.89530976374
			11'd1351: out = 32'b00000000000000001111001010111011; // input=-0.31982421875, output=1.89634028265
			11'd1352: out = 32'b00000000000000001111001011011101; // input=-0.32080078125, output=1.89737116015
			11'd1353: out = 32'b00000000000000001111001011111111; // input=-0.32177734375, output=1.89840239771
			11'd1354: out = 32'b00000000000000001111001100100001; // input=-0.32275390625, output=1.89943399682
			11'd1355: out = 32'b00000000000000001111001101000010; // input=-0.32373046875, output=1.90046595895
			11'd1356: out = 32'b00000000000000001111001101100100; // input=-0.32470703125, output=1.90149828559
			11'd1357: out = 32'b00000000000000001111001110000110; // input=-0.32568359375, output=1.90253097822
			11'd1358: out = 32'b00000000000000001111001110101000; // input=-0.32666015625, output=1.90356403834
			11'd1359: out = 32'b00000000000000001111001111001010; // input=-0.32763671875, output=1.90459746744
			11'd1360: out = 32'b00000000000000001111001111101100; // input=-0.32861328125, output=1.90563126703
			11'd1361: out = 32'b00000000000000001111010000001110; // input=-0.32958984375, output=1.9066654386
			11'd1362: out = 32'b00000000000000001111010000110000; // input=-0.33056640625, output=1.90769998367
			11'd1363: out = 32'b00000000000000001111010001010001; // input=-0.33154296875, output=1.90873490375
			11'd1364: out = 32'b00000000000000001111010001110011; // input=-0.33251953125, output=1.90977020035
			11'd1365: out = 32'b00000000000000001111010010010101; // input=-0.33349609375, output=1.91080587501
			11'd1366: out = 32'b00000000000000001111010010110111; // input=-0.33447265625, output=1.91184192924
			11'd1367: out = 32'b00000000000000001111010011011001; // input=-0.33544921875, output=1.91287836459
			11'd1368: out = 32'b00000000000000001111010011111011; // input=-0.33642578125, output=1.91391518257
			11'd1369: out = 32'b00000000000000001111010100011101; // input=-0.33740234375, output=1.91495238474
			11'd1370: out = 32'b00000000000000001111010100111111; // input=-0.33837890625, output=1.91598997263
			11'd1371: out = 32'b00000000000000001111010101100001; // input=-0.33935546875, output=1.9170279478
			11'd1372: out = 32'b00000000000000001111010110000011; // input=-0.34033203125, output=1.91806631181
			11'd1373: out = 32'b00000000000000001111010110100101; // input=-0.34130859375, output=1.9191050662
			11'd1374: out = 32'b00000000000000001111010111000111; // input=-0.34228515625, output=1.92014421254
			11'd1375: out = 32'b00000000000000001111010111101001; // input=-0.34326171875, output=1.9211837524
			11'd1376: out = 32'b00000000000000001111011000001011; // input=-0.34423828125, output=1.92222368735
			11'd1377: out = 32'b00000000000000001111011000101110; // input=-0.34521484375, output=1.92326401896
			11'd1378: out = 32'b00000000000000001111011001010000; // input=-0.34619140625, output=1.92430474883
			11'd1379: out = 32'b00000000000000001111011001110010; // input=-0.34716796875, output=1.92534587853
			11'd1380: out = 32'b00000000000000001111011010010100; // input=-0.34814453125, output=1.92638740965
			11'd1381: out = 32'b00000000000000001111011010110110; // input=-0.34912109375, output=1.9274293438
			11'd1382: out = 32'b00000000000000001111011011011000; // input=-0.35009765625, output=1.92847168257
			11'd1383: out = 32'b00000000000000001111011011111010; // input=-0.35107421875, output=1.92951442757
			11'd1384: out = 32'b00000000000000001111011100011101; // input=-0.35205078125, output=1.93055758041
			11'd1385: out = 32'b00000000000000001111011100111111; // input=-0.35302734375, output=1.9316011427
			11'd1386: out = 32'b00000000000000001111011101100001; // input=-0.35400390625, output=1.93264511606
			11'd1387: out = 32'b00000000000000001111011110000011; // input=-0.35498046875, output=1.93368950212
			11'd1388: out = 32'b00000000000000001111011110100101; // input=-0.35595703125, output=1.93473430252
			11'd1389: out = 32'b00000000000000001111011111001000; // input=-0.35693359375, output=1.93577951888
			11'd1390: out = 32'b00000000000000001111011111101010; // input=-0.35791015625, output=1.93682515284
			11'd1391: out = 32'b00000000000000001111100000001100; // input=-0.35888671875, output=1.93787120606
			11'd1392: out = 32'b00000000000000001111100000101110; // input=-0.35986328125, output=1.93891768017
			11'd1393: out = 32'b00000000000000001111100001010001; // input=-0.36083984375, output=1.93996457685
			11'd1394: out = 32'b00000000000000001111100001110011; // input=-0.36181640625, output=1.94101189774
			11'd1395: out = 32'b00000000000000001111100010010101; // input=-0.36279296875, output=1.94205964452
			11'd1396: out = 32'b00000000000000001111100010111000; // input=-0.36376953125, output=1.94310781886
			11'd1397: out = 32'b00000000000000001111100011011010; // input=-0.36474609375, output=1.94415642243
			11'd1398: out = 32'b00000000000000001111100011111100; // input=-0.36572265625, output=1.94520545691
			11'd1399: out = 32'b00000000000000001111100100011111; // input=-0.36669921875, output=1.946254924
			11'd1400: out = 32'b00000000000000001111100101000001; // input=-0.36767578125, output=1.94730482538
			11'd1401: out = 32'b00000000000000001111100101100100; // input=-0.36865234375, output=1.94835516276
			11'd1402: out = 32'b00000000000000001111100110000110; // input=-0.36962890625, output=1.94940593784
			11'd1403: out = 32'b00000000000000001111100110101001; // input=-0.37060546875, output=1.95045715233
			11'd1404: out = 32'b00000000000000001111100111001011; // input=-0.37158203125, output=1.95150880793
			11'd1405: out = 32'b00000000000000001111100111101110; // input=-0.37255859375, output=1.95256090639
			11'd1406: out = 32'b00000000000000001111101000010000; // input=-0.37353515625, output=1.95361344941
			11'd1407: out = 32'b00000000000000001111101000110011; // input=-0.37451171875, output=1.95466643873
			11'd1408: out = 32'b00000000000000001111101001010101; // input=-0.37548828125, output=1.95571987608
			11'd1409: out = 32'b00000000000000001111101001111000; // input=-0.37646484375, output=1.95677376322
			11'd1410: out = 32'b00000000000000001111101010011010; // input=-0.37744140625, output=1.95782810189
			11'd1411: out = 32'b00000000000000001111101010111101; // input=-0.37841796875, output=1.95888289384
			11'd1412: out = 32'b00000000000000001111101011011111; // input=-0.37939453125, output=1.95993814083
			11'd1413: out = 32'b00000000000000001111101100000010; // input=-0.38037109375, output=1.96099384464
			11'd1414: out = 32'b00000000000000001111101100100100; // input=-0.38134765625, output=1.96205000703
			11'd1415: out = 32'b00000000000000001111101101000111; // input=-0.38232421875, output=1.96310662977
			11'd1416: out = 32'b00000000000000001111101101101010; // input=-0.38330078125, output=1.96416371466
			11'd1417: out = 32'b00000000000000001111101110001100; // input=-0.38427734375, output=1.96522126348
			11'd1418: out = 32'b00000000000000001111101110101111; // input=-0.38525390625, output=1.96627927804
			11'd1419: out = 32'b00000000000000001111101111010010; // input=-0.38623046875, output=1.96733776012
			11'd1420: out = 32'b00000000000000001111101111110100; // input=-0.38720703125, output=1.96839671154
			11'd1421: out = 32'b00000000000000001111110000010111; // input=-0.38818359375, output=1.96945613411
			11'd1422: out = 32'b00000000000000001111110000111010; // input=-0.38916015625, output=1.97051602965
			11'd1423: out = 32'b00000000000000001111110001011101; // input=-0.39013671875, output=1.9715764
			11'd1424: out = 32'b00000000000000001111110001111111; // input=-0.39111328125, output=1.97263724697
			11'd1425: out = 32'b00000000000000001111110010100010; // input=-0.39208984375, output=1.97369857241
			11'd1426: out = 32'b00000000000000001111110011000101; // input=-0.39306640625, output=1.97476037817
			11'd1427: out = 32'b00000000000000001111110011101000; // input=-0.39404296875, output=1.9758226661
			11'd1428: out = 32'b00000000000000001111110100001011; // input=-0.39501953125, output=1.97688543805
			11'd1429: out = 32'b00000000000000001111110100101101; // input=-0.39599609375, output=1.97794869588
			11'd1430: out = 32'b00000000000000001111110101010000; // input=-0.39697265625, output=1.97901244148
			11'd1431: out = 32'b00000000000000001111110101110011; // input=-0.39794921875, output=1.98007667672
			11'd1432: out = 32'b00000000000000001111110110010110; // input=-0.39892578125, output=1.98114140347
			11'd1433: out = 32'b00000000000000001111110110111001; // input=-0.39990234375, output=1.98220662364
			11'd1434: out = 32'b00000000000000001111110111011100; // input=-0.40087890625, output=1.98327233911
			11'd1435: out = 32'b00000000000000001111110111111111; // input=-0.40185546875, output=1.98433855179
			11'd1436: out = 32'b00000000000000001111111000100010; // input=-0.40283203125, output=1.9854052636
			11'd1437: out = 32'b00000000000000001111111001000101; // input=-0.40380859375, output=1.98647247644
			11'd1438: out = 32'b00000000000000001111111001101000; // input=-0.40478515625, output=1.98754019225
			11'd1439: out = 32'b00000000000000001111111010001011; // input=-0.40576171875, output=1.98860841295
			11'd1440: out = 32'b00000000000000001111111010101110; // input=-0.40673828125, output=1.98967714048
			11'd1441: out = 32'b00000000000000001111111011010001; // input=-0.40771484375, output=1.99074637679
			11'd1442: out = 32'b00000000000000001111111011110100; // input=-0.40869140625, output=1.99181612382
			11'd1443: out = 32'b00000000000000001111111100010111; // input=-0.40966796875, output=1.99288638354
			11'd1444: out = 32'b00000000000000001111111100111010; // input=-0.41064453125, output=1.99395715791
			11'd1445: out = 32'b00000000000000001111111101011101; // input=-0.41162109375, output=1.9950284489
			11'd1446: out = 32'b00000000000000001111111110000000; // input=-0.41259765625, output=1.9961002585
			11'd1447: out = 32'b00000000000000001111111110100011; // input=-0.41357421875, output=1.99717258869
			11'd1448: out = 32'b00000000000000001111111111000111; // input=-0.41455078125, output=1.99824544146
			11'd1449: out = 32'b00000000000000001111111111101010; // input=-0.41552734375, output=1.99931881882
			11'd1450: out = 32'b00000000000000010000000000001101; // input=-0.41650390625, output=2.00039272277
			11'd1451: out = 32'b00000000000000010000000000110000; // input=-0.41748046875, output=2.00146715533
			11'd1452: out = 32'b00000000000000010000000001010011; // input=-0.41845703125, output=2.00254211853
			11'd1453: out = 32'b00000000000000010000000001110111; // input=-0.41943359375, output=2.00361761439
			11'd1454: out = 32'b00000000000000010000000010011010; // input=-0.42041015625, output=2.00469364496
			11'd1455: out = 32'b00000000000000010000000010111101; // input=-0.42138671875, output=2.00577021228
			11'd1456: out = 32'b00000000000000010000000011100000; // input=-0.42236328125, output=2.0068473184
			11'd1457: out = 32'b00000000000000010000000100000100; // input=-0.42333984375, output=2.00792496538
			11'd1458: out = 32'b00000000000000010000000100100111; // input=-0.42431640625, output=2.0090031553
			11'd1459: out = 32'b00000000000000010000000101001010; // input=-0.42529296875, output=2.01008189023
			11'd1460: out = 32'b00000000000000010000000101101110; // input=-0.42626953125, output=2.01116117226
			11'd1461: out = 32'b00000000000000010000000110010001; // input=-0.42724609375, output=2.01224100347
			11'd1462: out = 32'b00000000000000010000000110110101; // input=-0.42822265625, output=2.01332138597
			11'd1463: out = 32'b00000000000000010000000111011000; // input=-0.42919921875, output=2.01440232187
			11'd1464: out = 32'b00000000000000010000000111111011; // input=-0.43017578125, output=2.01548381328
			11'd1465: out = 32'b00000000000000010000001000011111; // input=-0.43115234375, output=2.01656586232
			11'd1466: out = 32'b00000000000000010000001001000010; // input=-0.43212890625, output=2.01764847113
			11'd1467: out = 32'b00000000000000010000001001100110; // input=-0.43310546875, output=2.01873164186
			11'd1468: out = 32'b00000000000000010000001010001001; // input=-0.43408203125, output=2.01981537664
			11'd1469: out = 32'b00000000000000010000001010101101; // input=-0.43505859375, output=2.02089967763
			11'd1470: out = 32'b00000000000000010000001011010000; // input=-0.43603515625, output=2.02198454701
			11'd1471: out = 32'b00000000000000010000001011110100; // input=-0.43701171875, output=2.02306998694
			11'd1472: out = 32'b00000000000000010000001100011000; // input=-0.43798828125, output=2.0241559996
			11'd1473: out = 32'b00000000000000010000001100111011; // input=-0.43896484375, output=2.02524258719
			11'd1474: out = 32'b00000000000000010000001101011111; // input=-0.43994140625, output=2.02632975191
			11'd1475: out = 32'b00000000000000010000001110000010; // input=-0.44091796875, output=2.02741749596
			11'd1476: out = 32'b00000000000000010000001110100110; // input=-0.44189453125, output=2.02850582155
			11'd1477: out = 32'b00000000000000010000001111001010; // input=-0.44287109375, output=2.02959473092
			11'd1478: out = 32'b00000000000000010000001111101101; // input=-0.44384765625, output=2.0306842263
			11'd1479: out = 32'b00000000000000010000010000010001; // input=-0.44482421875, output=2.03177430993
			11'd1480: out = 32'b00000000000000010000010000110101; // input=-0.44580078125, output=2.03286498406
			11'd1481: out = 32'b00000000000000010000010001011001; // input=-0.44677734375, output=2.03395625095
			11'd1482: out = 32'b00000000000000010000010001111100; // input=-0.44775390625, output=2.03504811287
			11'd1483: out = 32'b00000000000000010000010010100000; // input=-0.44873046875, output=2.0361405721
			11'd1484: out = 32'b00000000000000010000010011000100; // input=-0.44970703125, output=2.03723363093
			11'd1485: out = 32'b00000000000000010000010011101000; // input=-0.45068359375, output=2.03832729165
			11'd1486: out = 32'b00000000000000010000010100001100; // input=-0.45166015625, output=2.03942155657
			11'd1487: out = 32'b00000000000000010000010100110000; // input=-0.45263671875, output=2.040516428
			11'd1488: out = 32'b00000000000000010000010101010100; // input=-0.45361328125, output=2.04161190827
			11'd1489: out = 32'b00000000000000010000010101110111; // input=-0.45458984375, output=2.0427079997
			11'd1490: out = 32'b00000000000000010000010110011011; // input=-0.45556640625, output=2.04380470466
			11'd1491: out = 32'b00000000000000010000010110111111; // input=-0.45654296875, output=2.04490202548
			11'd1492: out = 32'b00000000000000010000010111100011; // input=-0.45751953125, output=2.04599996453
			11'd1493: out = 32'b00000000000000010000011000000111; // input=-0.45849609375, output=2.04709852418
			11'd1494: out = 32'b00000000000000010000011000101011; // input=-0.45947265625, output=2.04819770681
			11'd1495: out = 32'b00000000000000010000011001001111; // input=-0.46044921875, output=2.04929751482
			11'd1496: out = 32'b00000000000000010000011001110011; // input=-0.46142578125, output=2.0503979506
			11'd1497: out = 32'b00000000000000010000011010011000; // input=-0.46240234375, output=2.05149901657
			11'd1498: out = 32'b00000000000000010000011010111100; // input=-0.46337890625, output=2.05260071515
			11'd1499: out = 32'b00000000000000010000011011100000; // input=-0.46435546875, output=2.05370304877
			11'd1500: out = 32'b00000000000000010000011100000100; // input=-0.46533203125, output=2.05480601986
			11'd1501: out = 32'b00000000000000010000011100101000; // input=-0.46630859375, output=2.05590963089
			11'd1502: out = 32'b00000000000000010000011101001100; // input=-0.46728515625, output=2.05701388431
			11'd1503: out = 32'b00000000000000010000011101110000; // input=-0.46826171875, output=2.05811878259
			11'd1504: out = 32'b00000000000000010000011110010101; // input=-0.46923828125, output=2.05922432822
			11'd1505: out = 32'b00000000000000010000011110111001; // input=-0.47021484375, output=2.0603305237
			11'd1506: out = 32'b00000000000000010000011111011101; // input=-0.47119140625, output=2.06143737151
			11'd1507: out = 32'b00000000000000010000100000000001; // input=-0.47216796875, output=2.06254487418
			11'd1508: out = 32'b00000000000000010000100000100110; // input=-0.47314453125, output=2.06365303424
			11'd1509: out = 32'b00000000000000010000100001001010; // input=-0.47412109375, output=2.06476185421
			11'd1510: out = 32'b00000000000000010000100001101110; // input=-0.47509765625, output=2.06587133664
			11'd1511: out = 32'b00000000000000010000100010010011; // input=-0.47607421875, output=2.06698148409
			11'd1512: out = 32'b00000000000000010000100010110111; // input=-0.47705078125, output=2.06809229913
			11'd1513: out = 32'b00000000000000010000100011011100; // input=-0.47802734375, output=2.06920378434
			11'd1514: out = 32'b00000000000000010000100100000000; // input=-0.47900390625, output=2.0703159423
			11'd1515: out = 32'b00000000000000010000100100100101; // input=-0.47998046875, output=2.07142877563
			11'd1516: out = 32'b00000000000000010000100101001001; // input=-0.48095703125, output=2.07254228692
			11'd1517: out = 32'b00000000000000010000100101101110; // input=-0.48193359375, output=2.07365647881
			11'd1518: out = 32'b00000000000000010000100110010010; // input=-0.48291015625, output=2.07477135392
			11'd1519: out = 32'b00000000000000010000100110110111; // input=-0.48388671875, output=2.07588691492
			11'd1520: out = 32'b00000000000000010000100111011011; // input=-0.48486328125, output=2.07700316444
			11'd1521: out = 32'b00000000000000010000101000000000; // input=-0.48583984375, output=2.07812010518
			11'd1522: out = 32'b00000000000000010000101000100100; // input=-0.48681640625, output=2.07923773979
			11'd1523: out = 32'b00000000000000010000101001001001; // input=-0.48779296875, output=2.08035607099
			11'd1524: out = 32'b00000000000000010000101001101110; // input=-0.48876953125, output=2.08147510147
			11'd1525: out = 32'b00000000000000010000101010010010; // input=-0.48974609375, output=2.08259483396
			11'd1526: out = 32'b00000000000000010000101010110111; // input=-0.49072265625, output=2.08371527118
			11'd1527: out = 32'b00000000000000010000101011011100; // input=-0.49169921875, output=2.08483641586
			11'd1528: out = 32'b00000000000000010000101100000001; // input=-0.49267578125, output=2.08595827078
			11'd1529: out = 32'b00000000000000010000101100100101; // input=-0.49365234375, output=2.08708083869
			11'd1530: out = 32'b00000000000000010000101101001010; // input=-0.49462890625, output=2.08820412237
			11'd1531: out = 32'b00000000000000010000101101101111; // input=-0.49560546875, output=2.08932812462
			11'd1532: out = 32'b00000000000000010000101110010100; // input=-0.49658203125, output=2.09045284823
			11'd1533: out = 32'b00000000000000010000101110111001; // input=-0.49755859375, output=2.09157829602
			11'd1534: out = 32'b00000000000000010000101111011110; // input=-0.49853515625, output=2.09270447082
			11'd1535: out = 32'b00000000000000010000110000000011; // input=-0.49951171875, output=2.09383137548
			11'd1536: out = 32'b00000000000000010000110000101000; // input=-0.50048828125, output=2.09495901284
			11'd1537: out = 32'b00000000000000010000110001001101; // input=-0.50146484375, output=2.09608738578
			11'd1538: out = 32'b00000000000000010000110001110010; // input=-0.50244140625, output=2.09721649718
			11'd1539: out = 32'b00000000000000010000110010010111; // input=-0.50341796875, output=2.09834634992
			11'd1540: out = 32'b00000000000000010000110010111100; // input=-0.50439453125, output=2.09947694693
			11'd1541: out = 32'b00000000000000010000110011100001; // input=-0.50537109375, output=2.10060829111
			11'd1542: out = 32'b00000000000000010000110100000110; // input=-0.50634765625, output=2.1017403854
			11'd1543: out = 32'b00000000000000010000110100101011; // input=-0.50732421875, output=2.10287323276
			11'd1544: out = 32'b00000000000000010000110101010000; // input=-0.50830078125, output=2.10400683614
			11'd1545: out = 32'b00000000000000010000110101110101; // input=-0.50927734375, output=2.10514119851
			11'd1546: out = 32'b00000000000000010000110110011010; // input=-0.51025390625, output=2.10627632287
			11'd1547: out = 32'b00000000000000010000110111000000; // input=-0.51123046875, output=2.10741221223
			11'd1548: out = 32'b00000000000000010000110111100101; // input=-0.51220703125, output=2.10854886959
			11'd1549: out = 32'b00000000000000010000111000001010; // input=-0.51318359375, output=2.10968629798
			11'd1550: out = 32'b00000000000000010000111000101111; // input=-0.51416015625, output=2.11082450046
			11'd1551: out = 32'b00000000000000010000111001010101; // input=-0.51513671875, output=2.11196348009
			11'd1552: out = 32'b00000000000000010000111001111010; // input=-0.51611328125, output=2.11310323994
			11'd1553: out = 32'b00000000000000010000111010100000; // input=-0.51708984375, output=2.11424378309
			11'd1554: out = 32'b00000000000000010000111011000101; // input=-0.51806640625, output=2.11538511266
			11'd1555: out = 32'b00000000000000010000111011101010; // input=-0.51904296875, output=2.11652723175
			11'd1556: out = 32'b00000000000000010000111100010000; // input=-0.52001953125, output=2.11767014351
			11'd1557: out = 32'b00000000000000010000111100110101; // input=-0.52099609375, output=2.11881385109
			11'd1558: out = 32'b00000000000000010000111101011011; // input=-0.52197265625, output=2.11995835764
			11'd1559: out = 32'b00000000000000010000111110000000; // input=-0.52294921875, output=2.12110366635
			11'd1560: out = 32'b00000000000000010000111110100110; // input=-0.52392578125, output=2.12224978041
			11'd1561: out = 32'b00000000000000010000111111001011; // input=-0.52490234375, output=2.12339670303
			11'd1562: out = 32'b00000000000000010000111111110001; // input=-0.52587890625, output=2.12454443744
			11'd1563: out = 32'b00000000000000010001000000010111; // input=-0.52685546875, output=2.12569298688
			11'd1564: out = 32'b00000000000000010001000000111100; // input=-0.52783203125, output=2.1268423546
			11'd1565: out = 32'b00000000000000010001000001100010; // input=-0.52880859375, output=2.12799254388
			11'd1566: out = 32'b00000000000000010001000010001000; // input=-0.52978515625, output=2.12914355801
			11'd1567: out = 32'b00000000000000010001000010101110; // input=-0.53076171875, output=2.13029540029
			11'd1568: out = 32'b00000000000000010001000011010011; // input=-0.53173828125, output=2.13144807404
			11'd1569: out = 32'b00000000000000010001000011111001; // input=-0.53271484375, output=2.13260158261
			11'd1570: out = 32'b00000000000000010001000100011111; // input=-0.53369140625, output=2.13375592934
			11'd1571: out = 32'b00000000000000010001000101000101; // input=-0.53466796875, output=2.13491111761
			11'd1572: out = 32'b00000000000000010001000101101011; // input=-0.53564453125, output=2.13606715081
			11'd1573: out = 32'b00000000000000010001000110010001; // input=-0.53662109375, output=2.13722403234
			11'd1574: out = 32'b00000000000000010001000110110110; // input=-0.53759765625, output=2.13838176562
			11'd1575: out = 32'b00000000000000010001000111011100; // input=-0.53857421875, output=2.1395403541
			11'd1576: out = 32'b00000000000000010001001000000010; // input=-0.53955078125, output=2.14069980123
			11'd1577: out = 32'b00000000000000010001001000101000; // input=-0.54052734375, output=2.14186011048
			11'd1578: out = 32'b00000000000000010001001001001111; // input=-0.54150390625, output=2.14302128534
			11'd1579: out = 32'b00000000000000010001001001110101; // input=-0.54248046875, output=2.14418332933
			11'd1580: out = 32'b00000000000000010001001010011011; // input=-0.54345703125, output=2.14534624597
			11'd1581: out = 32'b00000000000000010001001011000001; // input=-0.54443359375, output=2.14651003881
			11'd1582: out = 32'b00000000000000010001001011100111; // input=-0.54541015625, output=2.14767471141
			11'd1583: out = 32'b00000000000000010001001100001101; // input=-0.54638671875, output=2.14884026735
			11'd1584: out = 32'b00000000000000010001001100110011; // input=-0.54736328125, output=2.15000671023
			11'd1585: out = 32'b00000000000000010001001101011010; // input=-0.54833984375, output=2.15117404367
			11'd1586: out = 32'b00000000000000010001001110000000; // input=-0.54931640625, output=2.15234227131
			11'd1587: out = 32'b00000000000000010001001110100110; // input=-0.55029296875, output=2.1535113968
			11'd1588: out = 32'b00000000000000010001001111001101; // input=-0.55126953125, output=2.15468142383
			11'd1589: out = 32'b00000000000000010001001111110011; // input=-0.55224609375, output=2.15585235607
			11'd1590: out = 32'b00000000000000010001010000011001; // input=-0.55322265625, output=2.15702419726
			11'd1591: out = 32'b00000000000000010001010001000000; // input=-0.55419921875, output=2.15819695111
			11'd1592: out = 32'b00000000000000010001010001100110; // input=-0.55517578125, output=2.15937062138
			11'd1593: out = 32'b00000000000000010001010010001101; // input=-0.55615234375, output=2.16054521185
			11'd1594: out = 32'b00000000000000010001010010110011; // input=-0.55712890625, output=2.1617207263
			11'd1595: out = 32'b00000000000000010001010011011010; // input=-0.55810546875, output=2.16289716856
			11'd1596: out = 32'b00000000000000010001010100000000; // input=-0.55908203125, output=2.16407454244
			11'd1597: out = 32'b00000000000000010001010100100111; // input=-0.56005859375, output=2.16525285181
			11'd1598: out = 32'b00000000000000010001010101001110; // input=-0.56103515625, output=2.16643210053
			11'd1599: out = 32'b00000000000000010001010101110100; // input=-0.56201171875, output=2.16761229251
			11'd1600: out = 32'b00000000000000010001010110011011; // input=-0.56298828125, output=2.16879343165
			11'd1601: out = 32'b00000000000000010001010111000010; // input=-0.56396484375, output=2.1699755219
			11'd1602: out = 32'b00000000000000010001010111101001; // input=-0.56494140625, output=2.1711585672
			11'd1603: out = 32'b00000000000000010001011000001111; // input=-0.56591796875, output=2.17234257154
			11'd1604: out = 32'b00000000000000010001011000110110; // input=-0.56689453125, output=2.17352753892
			11'd1605: out = 32'b00000000000000010001011001011101; // input=-0.56787109375, output=2.17471347335
			11'd1606: out = 32'b00000000000000010001011010000100; // input=-0.56884765625, output=2.17590037889
			11'd1607: out = 32'b00000000000000010001011010101011; // input=-0.56982421875, output=2.1770882596
			11'd1608: out = 32'b00000000000000010001011011010010; // input=-0.57080078125, output=2.17827711957
			11'd1609: out = 32'b00000000000000010001011011111001; // input=-0.57177734375, output=2.1794669629
			11'd1610: out = 32'b00000000000000010001011100100000; // input=-0.57275390625, output=2.18065779373
			11'd1611: out = 32'b00000000000000010001011101000111; // input=-0.57373046875, output=2.18184961621
			11'd1612: out = 32'b00000000000000010001011101101110; // input=-0.57470703125, output=2.18304243453
			11'd1613: out = 32'b00000000000000010001011110010101; // input=-0.57568359375, output=2.18423625289
			11'd1614: out = 32'b00000000000000010001011110111100; // input=-0.57666015625, output=2.1854310755
			11'd1615: out = 32'b00000000000000010001011111100011; // input=-0.57763671875, output=2.18662690663
			11'd1616: out = 32'b00000000000000010001100000001011; // input=-0.57861328125, output=2.18782375054
			11'd1617: out = 32'b00000000000000010001100000110010; // input=-0.57958984375, output=2.18902161152
			11'd1618: out = 32'b00000000000000010001100001011001; // input=-0.58056640625, output=2.19022049391
			11'd1619: out = 32'b00000000000000010001100010000000; // input=-0.58154296875, output=2.19142040204
			11'd1620: out = 32'b00000000000000010001100010101000; // input=-0.58251953125, output=2.19262134028
			11'd1621: out = 32'b00000000000000010001100011001111; // input=-0.58349609375, output=2.19382331303
			11'd1622: out = 32'b00000000000000010001100011110111; // input=-0.58447265625, output=2.1950263247
			11'd1623: out = 32'b00000000000000010001100100011110; // input=-0.58544921875, output=2.19623037975
			11'd1624: out = 32'b00000000000000010001100101000110; // input=-0.58642578125, output=2.19743548264
			11'd1625: out = 32'b00000000000000010001100101101101; // input=-0.58740234375, output=2.19864163786
			11'd1626: out = 32'b00000000000000010001100110010101; // input=-0.58837890625, output=2.19984884994
			11'd1627: out = 32'b00000000000000010001100110111100; // input=-0.58935546875, output=2.20105712342
			11'd1628: out = 32'b00000000000000010001100111100100; // input=-0.59033203125, output=2.20226646288
			11'd1629: out = 32'b00000000000000010001101000001100; // input=-0.59130859375, output=2.20347687291
			11'd1630: out = 32'b00000000000000010001101000110011; // input=-0.59228515625, output=2.20468835815
			11'd1631: out = 32'b00000000000000010001101001011011; // input=-0.59326171875, output=2.20590092324
			11'd1632: out = 32'b00000000000000010001101010000011; // input=-0.59423828125, output=2.20711457287
			11'd1633: out = 32'b00000000000000010001101010101011; // input=-0.59521484375, output=2.20832931175
			11'd1634: out = 32'b00000000000000010001101011010010; // input=-0.59619140625, output=2.2095451446
			11'd1635: out = 32'b00000000000000010001101011111010; // input=-0.59716796875, output=2.21076207619
			11'd1636: out = 32'b00000000000000010001101100100010; // input=-0.59814453125, output=2.21198011132
			11'd1637: out = 32'b00000000000000010001101101001010; // input=-0.59912109375, output=2.21319925481
			11'd1638: out = 32'b00000000000000010001101101110010; // input=-0.60009765625, output=2.21441951149
			11'd1639: out = 32'b00000000000000010001101110011010; // input=-0.60107421875, output=2.21564088625
			11'd1640: out = 32'b00000000000000010001101111000010; // input=-0.60205078125, output=2.216863384
			11'd1641: out = 32'b00000000000000010001101111101010; // input=-0.60302734375, output=2.21808700967
			11'd1642: out = 32'b00000000000000010001110000010010; // input=-0.60400390625, output=2.21931176822
			11'd1643: out = 32'b00000000000000010001110000111011; // input=-0.60498046875, output=2.22053766465
			11'd1644: out = 32'b00000000000000010001110001100011; // input=-0.60595703125, output=2.22176470399
			11'd1645: out = 32'b00000000000000010001110010001011; // input=-0.60693359375, output=2.22299289128
			11'd1646: out = 32'b00000000000000010001110010110011; // input=-0.60791015625, output=2.22422223162
			11'd1647: out = 32'b00000000000000010001110011011100; // input=-0.60888671875, output=2.22545273013
			11'd1648: out = 32'b00000000000000010001110100000100; // input=-0.60986328125, output=2.22668439194
			11'd1649: out = 32'b00000000000000010001110100101100; // input=-0.61083984375, output=2.22791722224
			11'd1650: out = 32'b00000000000000010001110101010101; // input=-0.61181640625, output=2.22915122625
			11'd1651: out = 32'b00000000000000010001110101111101; // input=-0.61279296875, output=2.23038640919
			11'd1652: out = 32'b00000000000000010001110110100110; // input=-0.61376953125, output=2.23162277636
			11'd1653: out = 32'b00000000000000010001110111001110; // input=-0.61474609375, output=2.23286033305
			11'd1654: out = 32'b00000000000000010001110111110111; // input=-0.61572265625, output=2.23409908462
			11'd1655: out = 32'b00000000000000010001111000100000; // input=-0.61669921875, output=2.23533903642
			11'd1656: out = 32'b00000000000000010001111001001000; // input=-0.61767578125, output=2.23658019387
			11'd1657: out = 32'b00000000000000010001111001110001; // input=-0.61865234375, output=2.23782256242
			11'd1658: out = 32'b00000000000000010001111010011010; // input=-0.61962890625, output=2.23906614753
			11'd1659: out = 32'b00000000000000010001111011000011; // input=-0.62060546875, output=2.24031095471
			11'd1660: out = 32'b00000000000000010001111011101011; // input=-0.62158203125, output=2.24155698952
			11'd1661: out = 32'b00000000000000010001111100010100; // input=-0.62255859375, output=2.24280425753
			11'd1662: out = 32'b00000000000000010001111100111101; // input=-0.62353515625, output=2.24405276435
			11'd1663: out = 32'b00000000000000010001111101100110; // input=-0.62451171875, output=2.24530251564
			11'd1664: out = 32'b00000000000000010001111110001111; // input=-0.62548828125, output=2.24655351708
			11'd1665: out = 32'b00000000000000010001111110111000; // input=-0.62646484375, output=2.24780577439
			11'd1666: out = 32'b00000000000000010001111111100001; // input=-0.62744140625, output=2.24905929334
			11'd1667: out = 32'b00000000000000010010000000001010; // input=-0.62841796875, output=2.25031407972
			11'd1668: out = 32'b00000000000000010010000000110011; // input=-0.62939453125, output=2.25157013937
			11'd1669: out = 32'b00000000000000010010000001011101; // input=-0.63037109375, output=2.25282747815
			11'd1670: out = 32'b00000000000000010010000010000110; // input=-0.63134765625, output=2.25408610198
			11'd1671: out = 32'b00000000000000010010000010101111; // input=-0.63232421875, output=2.25534601681
			11'd1672: out = 32'b00000000000000010010000011011001; // input=-0.63330078125, output=2.25660722861
			11'd1673: out = 32'b00000000000000010010000100000010; // input=-0.63427734375, output=2.25786974343
			11'd1674: out = 32'b00000000000000010010000100101011; // input=-0.63525390625, output=2.25913356731
			11'd1675: out = 32'b00000000000000010010000101010101; // input=-0.63623046875, output=2.26039870638
			11'd1676: out = 32'b00000000000000010010000101111110; // input=-0.63720703125, output=2.26166516677
			11'd1677: out = 32'b00000000000000010010000110101000; // input=-0.63818359375, output=2.26293295467
			11'd1678: out = 32'b00000000000000010010000111010001; // input=-0.63916015625, output=2.26420207631
			11'd1679: out = 32'b00000000000000010010000111111011; // input=-0.64013671875, output=2.26547253796
			11'd1680: out = 32'b00000000000000010010001000100101; // input=-0.64111328125, output=2.26674434592
			11'd1681: out = 32'b00000000000000010010001001001110; // input=-0.64208984375, output=2.26801750655
			11'd1682: out = 32'b00000000000000010010001001111000; // input=-0.64306640625, output=2.26929202626
			11'd1683: out = 32'b00000000000000010010001010100010; // input=-0.64404296875, output=2.27056791146
			11'd1684: out = 32'b00000000000000010010001011001100; // input=-0.64501953125, output=2.27184516865
			11'd1685: out = 32'b00000000000000010010001011110110; // input=-0.64599609375, output=2.27312380436
			11'd1686: out = 32'b00000000000000010010001100100000; // input=-0.64697265625, output=2.27440382515
			11'd1687: out = 32'b00000000000000010010001101001010; // input=-0.64794921875, output=2.27568523764
			11'd1688: out = 32'b00000000000000010010001101110100; // input=-0.64892578125, output=2.27696804848
			11'd1689: out = 32'b00000000000000010010001110011110; // input=-0.64990234375, output=2.27825226439
			11'd1690: out = 32'b00000000000000010010001111001000; // input=-0.65087890625, output=2.27953789212
			11'd1691: out = 32'b00000000000000010010001111110010; // input=-0.65185546875, output=2.28082493846
			11'd1692: out = 32'b00000000000000010010010000011100; // input=-0.65283203125, output=2.28211341026
			11'd1693: out = 32'b00000000000000010010010001000111; // input=-0.65380859375, output=2.28340331442
			11'd1694: out = 32'b00000000000000010010010001110001; // input=-0.65478515625, output=2.28469465787
			11'd1695: out = 32'b00000000000000010010010010011011; // input=-0.65576171875, output=2.2859874476
			11'd1696: out = 32'b00000000000000010010010011000110; // input=-0.65673828125, output=2.28728169065
			11'd1697: out = 32'b00000000000000010010010011110000; // input=-0.65771484375, output=2.28857739412
			11'd1698: out = 32'b00000000000000010010010100011011; // input=-0.65869140625, output=2.28987456513
			11'd1699: out = 32'b00000000000000010010010101000101; // input=-0.65966796875, output=2.29117321088
			11'd1700: out = 32'b00000000000000010010010101110000; // input=-0.66064453125, output=2.2924733386
			11'd1701: out = 32'b00000000000000010010010110011010; // input=-0.66162109375, output=2.29377495559
			11'd1702: out = 32'b00000000000000010010010111000101; // input=-0.66259765625, output=2.29507806919
			11'd1703: out = 32'b00000000000000010010010111110000; // input=-0.66357421875, output=2.29638268678
			11'd1704: out = 32'b00000000000000010010011000011011; // input=-0.66455078125, output=2.29768881583
			11'd1705: out = 32'b00000000000000010010011001000110; // input=-0.66552734375, output=2.29899646382
			11'd1706: out = 32'b00000000000000010010011001110000; // input=-0.66650390625, output=2.30030563833
			11'd1707: out = 32'b00000000000000010010011010011011; // input=-0.66748046875, output=2.30161634695
			11'd1708: out = 32'b00000000000000010010011011000110; // input=-0.66845703125, output=2.30292859735
			11'd1709: out = 32'b00000000000000010010011011110001; // input=-0.66943359375, output=2.30424239726
			11'd1710: out = 32'b00000000000000010010011100011101; // input=-0.67041015625, output=2.30555775445
			11'd1711: out = 32'b00000000000000010010011101001000; // input=-0.67138671875, output=2.30687467675
			11'd1712: out = 32'b00000000000000010010011101110011; // input=-0.67236328125, output=2.30819317206
			11'd1713: out = 32'b00000000000000010010011110011110; // input=-0.67333984375, output=2.30951324833
			11'd1714: out = 32'b00000000000000010010011111001001; // input=-0.67431640625, output=2.31083491357
			11'd1715: out = 32'b00000000000000010010011111110101; // input=-0.67529296875, output=2.31215817585
			11'd1716: out = 32'b00000000000000010010100000100000; // input=-0.67626953125, output=2.3134830433
			11'd1717: out = 32'b00000000000000010010100001001100; // input=-0.67724609375, output=2.3148095241
			11'd1718: out = 32'b00000000000000010010100001110111; // input=-0.67822265625, output=2.3161376265
			11'd1719: out = 32'b00000000000000010010100010100011; // input=-0.67919921875, output=2.31746735883
			11'd1720: out = 32'b00000000000000010010100011001110; // input=-0.68017578125, output=2.31879872945
			11'd1721: out = 32'b00000000000000010010100011111010; // input=-0.68115234375, output=2.32013174681
			11'd1722: out = 32'b00000000000000010010100100100110; // input=-0.68212890625, output=2.3214664194
			11'd1723: out = 32'b00000000000000010010100101010010; // input=-0.68310546875, output=2.3228027558
			11'd1724: out = 32'b00000000000000010010100101111101; // input=-0.68408203125, output=2.32414076463
			11'd1725: out = 32'b00000000000000010010100110101001; // input=-0.68505859375, output=2.32548045461
			11'd1726: out = 32'b00000000000000010010100111010101; // input=-0.68603515625, output=2.32682183449
			11'd1727: out = 32'b00000000000000010010101000000001; // input=-0.68701171875, output=2.32816491311
			11'd1728: out = 32'b00000000000000010010101000101101; // input=-0.68798828125, output=2.32950969936
			11'd1729: out = 32'b00000000000000010010101001011001; // input=-0.68896484375, output=2.33085620223
			11'd1730: out = 32'b00000000000000010010101010000110; // input=-0.68994140625, output=2.33220443076
			11'd1731: out = 32'b00000000000000010010101010110010; // input=-0.69091796875, output=2.33355439404
			11'd1732: out = 32'b00000000000000010010101011011110; // input=-0.69189453125, output=2.33490610128
			11'd1733: out = 32'b00000000000000010010101100001011; // input=-0.69287109375, output=2.33625956172
			11'd1734: out = 32'b00000000000000010010101100110111; // input=-0.69384765625, output=2.33761478469
			11'd1735: out = 32'b00000000000000010010101101100011; // input=-0.69482421875, output=2.3389717796
			11'd1736: out = 32'b00000000000000010010101110010000; // input=-0.69580078125, output=2.34033055592
			11'd1737: out = 32'b00000000000000010010101110111101; // input=-0.69677734375, output=2.34169112321
			11'd1738: out = 32'b00000000000000010010101111101001; // input=-0.69775390625, output=2.34305349109
			11'd1739: out = 32'b00000000000000010010110000010110; // input=-0.69873046875, output=2.34441766927
			11'd1740: out = 32'b00000000000000010010110001000011; // input=-0.69970703125, output=2.34578366754
			11'd1741: out = 32'b00000000000000010010110001101111; // input=-0.70068359375, output=2.34715149575
			11'd1742: out = 32'b00000000000000010010110010011100; // input=-0.70166015625, output=2.34852116386
			11'd1743: out = 32'b00000000000000010010110011001001; // input=-0.70263671875, output=2.34989268189
			11'd1744: out = 32'b00000000000000010010110011110110; // input=-0.70361328125, output=2.35126605994
			11'd1745: out = 32'b00000000000000010010110100100011; // input=-0.70458984375, output=2.3526413082
			11'd1746: out = 32'b00000000000000010010110101010000; // input=-0.70556640625, output=2.35401843695
			11'd1747: out = 32'b00000000000000010010110101111110; // input=-0.70654296875, output=2.35539745654
			11'd1748: out = 32'b00000000000000010010110110101011; // input=-0.70751953125, output=2.35677837743
			11'd1749: out = 32'b00000000000000010010110111011000; // input=-0.70849609375, output=2.35816121012
			11'd1750: out = 32'b00000000000000010010111000000110; // input=-0.70947265625, output=2.35954596526
			11'd1751: out = 32'b00000000000000010010111000110011; // input=-0.71044921875, output=2.36093265353
			11'd1752: out = 32'b00000000000000010010111001100001; // input=-0.71142578125, output=2.36232128574
			11'd1753: out = 32'b00000000000000010010111010001110; // input=-0.71240234375, output=2.36371187278
			11'd1754: out = 32'b00000000000000010010111010111100; // input=-0.71337890625, output=2.36510442562
			11'd1755: out = 32'b00000000000000010010111011101001; // input=-0.71435546875, output=2.36649895534
			11'd1756: out = 32'b00000000000000010010111100010111; // input=-0.71533203125, output=2.36789547311
			11'd1757: out = 32'b00000000000000010010111101000101; // input=-0.71630859375, output=2.36929399018
			11'd1758: out = 32'b00000000000000010010111101110011; // input=-0.71728515625, output=2.37069451791
			11'd1759: out = 32'b00000000000000010010111110100001; // input=-0.71826171875, output=2.37209706777
			11'd1760: out = 32'b00000000000000010010111111001111; // input=-0.71923828125, output=2.3735016513
			11'd1761: out = 32'b00000000000000010010111111111101; // input=-0.72021484375, output=2.37490828016
			11'd1762: out = 32'b00000000000000010011000000101011; // input=-0.72119140625, output=2.37631696612
			11'd1763: out = 32'b00000000000000010011000001011001; // input=-0.72216796875, output=2.37772772102
			11'd1764: out = 32'b00000000000000010011000010001000; // input=-0.72314453125, output=2.37914055683
			11'd1765: out = 32'b00000000000000010011000010110110; // input=-0.72412109375, output=2.38055548562
			11'd1766: out = 32'b00000000000000010011000011100100; // input=-0.72509765625, output=2.38197251956
			11'd1767: out = 32'b00000000000000010011000100010011; // input=-0.72607421875, output=2.38339167094
			11'd1768: out = 32'b00000000000000010011000101000010; // input=-0.72705078125, output=2.38481295214
			11'd1769: out = 32'b00000000000000010011000101110000; // input=-0.72802734375, output=2.38623637568
			11'd1770: out = 32'b00000000000000010011000110011111; // input=-0.72900390625, output=2.38766195416
			11'd1771: out = 32'b00000000000000010011000111001110; // input=-0.72998046875, output=2.38908970031
			11'd1772: out = 32'b00000000000000010011000111111101; // input=-0.73095703125, output=2.39051962697
			11'd1773: out = 32'b00000000000000010011001000101011; // input=-0.73193359375, output=2.3919517471
			11'd1774: out = 32'b00000000000000010011001001011010; // input=-0.73291015625, output=2.39338607378
			11'd1775: out = 32'b00000000000000010011001010001010; // input=-0.73388671875, output=2.39482262021
			11'd1776: out = 32'b00000000000000010011001010111001; // input=-0.73486328125, output=2.39626139969
			11'd1777: out = 32'b00000000000000010011001011101000; // input=-0.73583984375, output=2.39770242567
			11'd1778: out = 32'b00000000000000010011001100010111; // input=-0.73681640625, output=2.39914571171
			11'd1779: out = 32'b00000000000000010011001101000111; // input=-0.73779296875, output=2.4005912715
			11'd1780: out = 32'b00000000000000010011001101110110; // input=-0.73876953125, output=2.40203911885
			11'd1781: out = 32'b00000000000000010011001110100110; // input=-0.73974609375, output=2.40348926771
			11'd1782: out = 32'b00000000000000010011001111010101; // input=-0.74072265625, output=2.40494173215
			11'd1783: out = 32'b00000000000000010011010000000101; // input=-0.74169921875, output=2.40639652638
			11'd1784: out = 32'b00000000000000010011010000110101; // input=-0.74267578125, output=2.40785366474
			11'd1785: out = 32'b00000000000000010011010001100100; // input=-0.74365234375, output=2.40931316171
			11'd1786: out = 32'b00000000000000010011010010010100; // input=-0.74462890625, output=2.4107750319
			11'd1787: out = 32'b00000000000000010011010011000100; // input=-0.74560546875, output=2.41223929006
			11'd1788: out = 32'b00000000000000010011010011110100; // input=-0.74658203125, output=2.4137059511
			11'd1789: out = 32'b00000000000000010011010100100100; // input=-0.74755859375, output=2.41517503004
			11'd1790: out = 32'b00000000000000010011010101010101; // input=-0.74853515625, output=2.41664654208
			11'd1791: out = 32'b00000000000000010011010110000101; // input=-0.74951171875, output=2.41812050255
			11'd1792: out = 32'b00000000000000010011010110110101; // input=-0.75048828125, output=2.41959692693
			11'd1793: out = 32'b00000000000000010011010111100110; // input=-0.75146484375, output=2.42107583084
			11'd1794: out = 32'b00000000000000010011011000010110; // input=-0.75244140625, output=2.42255723008
			11'd1795: out = 32'b00000000000000010011011001000111; // input=-0.75341796875, output=2.42404114058
			11'd1796: out = 32'b00000000000000010011011001111000; // input=-0.75439453125, output=2.42552757845
			11'd1797: out = 32'b00000000000000010011011010101000; // input=-0.75537109375, output=2.42701655995
			11'd1798: out = 32'b00000000000000010011011011011001; // input=-0.75634765625, output=2.42850810149
			11'd1799: out = 32'b00000000000000010011011100001010; // input=-0.75732421875, output=2.43000221966
			11'd1800: out = 32'b00000000000000010011011100111011; // input=-0.75830078125, output=2.43149893121
			11'd1801: out = 32'b00000000000000010011011101101100; // input=-0.75927734375, output=2.43299825307
			11'd1802: out = 32'b00000000000000010011011110011110; // input=-0.76025390625, output=2.43450020233
			11'd1803: out = 32'b00000000000000010011011111001111; // input=-0.76123046875, output=2.43600479626
			11'd1804: out = 32'b00000000000000010011100000000000; // input=-0.76220703125, output=2.4375120523
			11'd1805: out = 32'b00000000000000010011100000110010; // input=-0.76318359375, output=2.43902198807
			11'd1806: out = 32'b00000000000000010011100001100011; // input=-0.76416015625, output=2.44053462137
			11'd1807: out = 32'b00000000000000010011100010010101; // input=-0.76513671875, output=2.44204997021
			11'd1808: out = 32'b00000000000000010011100011000111; // input=-0.76611328125, output=2.44356805275
			11'd1809: out = 32'b00000000000000010011100011111001; // input=-0.76708984375, output=2.44508888736
			11'd1810: out = 32'b00000000000000010011100100101011; // input=-0.76806640625, output=2.44661249259
			11'd1811: out = 32'b00000000000000010011100101011101; // input=-0.76904296875, output=2.44813888721
			11'd1812: out = 32'b00000000000000010011100110001111; // input=-0.77001953125, output=2.44966809017
			11'd1813: out = 32'b00000000000000010011100111000001; // input=-0.77099609375, output=2.45120012061
			11'd1814: out = 32'b00000000000000010011100111110011; // input=-0.77197265625, output=2.4527349979
			11'd1815: out = 32'b00000000000000010011101000100110; // input=-0.77294921875, output=2.45427274161
			11'd1816: out = 32'b00000000000000010011101001011000; // input=-0.77392578125, output=2.4558133715
			11'd1817: out = 32'b00000000000000010011101010001011; // input=-0.77490234375, output=2.45735690757
			11'd1818: out = 32'b00000000000000010011101010111101; // input=-0.77587890625, output=2.45890337003
			11'd1819: out = 32'b00000000000000010011101011110000; // input=-0.77685546875, output=2.4604527793
			11'd1820: out = 32'b00000000000000010011101100100011; // input=-0.77783203125, output=2.46200515604
			11'd1821: out = 32'b00000000000000010011101101010110; // input=-0.77880859375, output=2.46356052112
			11'd1822: out = 32'b00000000000000010011101110001001; // input=-0.77978515625, output=2.46511889565
			11'd1823: out = 32'b00000000000000010011101110111100; // input=-0.78076171875, output=2.46668030098
			11'd1824: out = 32'b00000000000000010011101111101111; // input=-0.78173828125, output=2.46824475868
			11'd1825: out = 32'b00000000000000010011110000100011; // input=-0.78271484375, output=2.46981229058
			11'd1826: out = 32'b00000000000000010011110001010110; // input=-0.78369140625, output=2.47138291876
			11'd1827: out = 32'b00000000000000010011110010001010; // input=-0.78466796875, output=2.47295666552
			11'd1828: out = 32'b00000000000000010011110010111110; // input=-0.78564453125, output=2.47453355344
			11'd1829: out = 32'b00000000000000010011110011110001; // input=-0.78662109375, output=2.47611360534
			11'd1830: out = 32'b00000000000000010011110100100101; // input=-0.78759765625, output=2.47769684433
			11'd1831: out = 32'b00000000000000010011110101011001; // input=-0.78857421875, output=2.47928329375
			11'd1832: out = 32'b00000000000000010011110110001101; // input=-0.78955078125, output=2.48087297723
			11'd1833: out = 32'b00000000000000010011110111000001; // input=-0.79052734375, output=2.48246591868
			11'd1834: out = 32'b00000000000000010011110111110110; // input=-0.79150390625, output=2.48406214227
			11'd1835: out = 32'b00000000000000010011111000101010; // input=-0.79248046875, output=2.48566167247
			11'd1836: out = 32'b00000000000000010011111001011111; // input=-0.79345703125, output=2.48726453403
			11'd1837: out = 32'b00000000000000010011111010010011; // input=-0.79443359375, output=2.488870752
			11'd1838: out = 32'b00000000000000010011111011001000; // input=-0.79541015625, output=2.49048035171
			11'd1839: out = 32'b00000000000000010011111011111101; // input=-0.79638671875, output=2.49209335883
			11'd1840: out = 32'b00000000000000010011111100110010; // input=-0.79736328125, output=2.4937097993
			11'd1841: out = 32'b00000000000000010011111101100111; // input=-0.79833984375, output=2.49532969939
			11'd1842: out = 32'b00000000000000010011111110011100; // input=-0.79931640625, output=2.49695308569
			11'd1843: out = 32'b00000000000000010011111111010001; // input=-0.80029296875, output=2.49857998512
			11'd1844: out = 32'b00000000000000010100000000000111; // input=-0.80126953125, output=2.5002104249
			11'd1845: out = 32'b00000000000000010100000000111100; // input=-0.80224609375, output=2.50184443262
			11'd1846: out = 32'b00000000000000010100000001110010; // input=-0.80322265625, output=2.5034820362
			11'd1847: out = 32'b00000000000000010100000010101000; // input=-0.80419921875, output=2.50512326391
			11'd1848: out = 32'b00000000000000010100000011011110; // input=-0.80517578125, output=2.50676814435
			11'd1849: out = 32'b00000000000000010100000100010100; // input=-0.80615234375, output=2.50841670652
			11'd1850: out = 32'b00000000000000010100000101001010; // input=-0.80712890625, output=2.51006897974
			11'd1851: out = 32'b00000000000000010100000110000000; // input=-0.80810546875, output=2.51172499375
			11'd1852: out = 32'b00000000000000010100000110110111; // input=-0.80908203125, output=2.51338477864
			11'd1853: out = 32'b00000000000000010100000111101101; // input=-0.81005859375, output=2.51504836488
			11'd1854: out = 32'b00000000000000010100001000100100; // input=-0.81103515625, output=2.51671578336
			11'd1855: out = 32'b00000000000000010100001001011011; // input=-0.81201171875, output=2.51838706534
			11'd1856: out = 32'b00000000000000010100001010010001; // input=-0.81298828125, output=2.52006224252
			11'd1857: out = 32'b00000000000000010100001011001000; // input=-0.81396484375, output=2.52174134698
			11'd1858: out = 32'b00000000000000010100001100000000; // input=-0.81494140625, output=2.52342441124
			11'd1859: out = 32'b00000000000000010100001100110111; // input=-0.81591796875, output=2.52511146826
			11'd1860: out = 32'b00000000000000010100001101101110; // input=-0.81689453125, output=2.52680255142
			11'd1861: out = 32'b00000000000000010100001110100110; // input=-0.81787109375, output=2.52849769456
			11'd1862: out = 32'b00000000000000010100001111011101; // input=-0.81884765625, output=2.53019693197
			11'd1863: out = 32'b00000000000000010100010000010101; // input=-0.81982421875, output=2.53190029839
			11'd1864: out = 32'b00000000000000010100010001001101; // input=-0.82080078125, output=2.53360782906
			11'd1865: out = 32'b00000000000000010100010010000101; // input=-0.82177734375, output=2.53531955968
			11'd1866: out = 32'b00000000000000010100010010111110; // input=-0.82275390625, output=2.53703552645
			11'd1867: out = 32'b00000000000000010100010011110110; // input=-0.82373046875, output=2.53875576607
			11'd1868: out = 32'b00000000000000010100010100101110; // input=-0.82470703125, output=2.54048031574
			11'd1869: out = 32'b00000000000000010100010101100111; // input=-0.82568359375, output=2.54220921319
			11'd1870: out = 32'b00000000000000010100010110100000; // input=-0.82666015625, output=2.54394249668
			11'd1871: out = 32'b00000000000000010100010111011001; // input=-0.82763671875, output=2.54568020501
			11'd1872: out = 32'b00000000000000010100011000010010; // input=-0.82861328125, output=2.54742237753
			11'd1873: out = 32'b00000000000000010100011001001011; // input=-0.82958984375, output=2.54916905414
			11'd1874: out = 32'b00000000000000010100011010000101; // input=-0.83056640625, output=2.55092027535
			11'd1875: out = 32'b00000000000000010100011010111110; // input=-0.83154296875, output=2.55267608221
			11'd1876: out = 32'b00000000000000010100011011111000; // input=-0.83251953125, output=2.5544365164
			11'd1877: out = 32'b00000000000000010100011100110010; // input=-0.83349609375, output=2.55620162019
			11'd1878: out = 32'b00000000000000010100011101101100; // input=-0.83447265625, output=2.55797143649
			11'd1879: out = 32'b00000000000000010100011110100110; // input=-0.83544921875, output=2.55974600883
			11'd1880: out = 32'b00000000000000010100011111100000; // input=-0.83642578125, output=2.5615253814
			11'd1881: out = 32'b00000000000000010100100000011011; // input=-0.83740234375, output=2.56330959903
			11'd1882: out = 32'b00000000000000010100100001010101; // input=-0.83837890625, output=2.56509870727
			11'd1883: out = 32'b00000000000000010100100010010000; // input=-0.83935546875, output=2.5668927523
			11'd1884: out = 32'b00000000000000010100100011001011; // input=-0.84033203125, output=2.56869178106
			11'd1885: out = 32'b00000000000000010100100100000110; // input=-0.84130859375, output=2.57049584118
			11'd1886: out = 32'b00000000000000010100100101000001; // input=-0.84228515625, output=2.57230498103
			11'd1887: out = 32'b00000000000000010100100101111101; // input=-0.84326171875, output=2.57411924973
			11'd1888: out = 32'b00000000000000010100100110111000; // input=-0.84423828125, output=2.57593869719
			11'd1889: out = 32'b00000000000000010100100111110100; // input=-0.84521484375, output=2.57776337407
			11'd1890: out = 32'b00000000000000010100101000110000; // input=-0.84619140625, output=2.57959333186
			11'd1891: out = 32'b00000000000000010100101001101100; // input=-0.84716796875, output=2.58142862285
			11'd1892: out = 32'b00000000000000010100101010101001; // input=-0.84814453125, output=2.58326930019
			11'd1893: out = 32'b00000000000000010100101011100101; // input=-0.84912109375, output=2.58511541787
			11'd1894: out = 32'b00000000000000010100101100100010; // input=-0.85009765625, output=2.58696703077
			11'd1895: out = 32'b00000000000000010100101101011111; // input=-0.85107421875, output=2.58882419465
			11'd1896: out = 32'b00000000000000010100101110011100; // input=-0.85205078125, output=2.59068696621
			11'd1897: out = 32'b00000000000000010100101111011001; // input=-0.85302734375, output=2.59255540308
			11'd1898: out = 32'b00000000000000010100110000010110; // input=-0.85400390625, output=2.59442956385
			11'd1899: out = 32'b00000000000000010100110001010100; // input=-0.85498046875, output=2.59630950808
			11'd1900: out = 32'b00000000000000010100110010010010; // input=-0.85595703125, output=2.59819529636
			11'd1901: out = 32'b00000000000000010100110011010000; // input=-0.85693359375, output=2.60008699031
			11'd1902: out = 32'b00000000000000010100110100001110; // input=-0.85791015625, output=2.60198465258
			11'd1903: out = 32'b00000000000000010100110101001100; // input=-0.85888671875, output=2.60388834693
			11'd1904: out = 32'b00000000000000010100110110001011; // input=-0.85986328125, output=2.60579813822
			11'd1905: out = 32'b00000000000000010100110111001010; // input=-0.86083984375, output=2.60771409243
			11'd1906: out = 32'b00000000000000010100111000001001; // input=-0.86181640625, output=2.60963627672
			11'd1907: out = 32'b00000000000000010100111001001000; // input=-0.86279296875, output=2.61156475943
			11'd1908: out = 32'b00000000000000010100111010000111; // input=-0.86376953125, output=2.61349961013
			11'd1909: out = 32'b00000000000000010100111011000111; // input=-0.86474609375, output=2.61544089964
			11'd1910: out = 32'b00000000000000010100111100000111; // input=-0.86572265625, output=2.61738870006
			11'd1911: out = 32'b00000000000000010100111101000111; // input=-0.86669921875, output=2.61934308481
			11'd1912: out = 32'b00000000000000010100111110000111; // input=-0.86767578125, output=2.62130412866
			11'd1913: out = 32'b00000000000000010100111111000111; // input=-0.86865234375, output=2.62327190776
			11'd1914: out = 32'b00000000000000010101000000001000; // input=-0.86962890625, output=2.62524649969
			11'd1915: out = 32'b00000000000000010101000001001001; // input=-0.87060546875, output=2.62722798349
			11'd1916: out = 32'b00000000000000010101000010001010; // input=-0.87158203125, output=2.62921643969
			11'd1917: out = 32'b00000000000000010101000011001100; // input=-0.87255859375, output=2.63121195036
			11'd1918: out = 32'b00000000000000010101000100001101; // input=-0.87353515625, output=2.63321459915
			11'd1919: out = 32'b00000000000000010101000101001111; // input=-0.87451171875, output=2.63522447134
			11'd1920: out = 32'b00000000000000010101000110010001; // input=-0.87548828125, output=2.63724165386
			11'd1921: out = 32'b00000000000000010101000111010011; // input=-0.87646484375, output=2.63926623536
			11'd1922: out = 32'b00000000000000010101001000010110; // input=-0.87744140625, output=2.64129830626
			11'd1923: out = 32'b00000000000000010101001001011001; // input=-0.87841796875, output=2.64333795878
			11'd1924: out = 32'b00000000000000010101001010011100; // input=-0.87939453125, output=2.645385287
			11'd1925: out = 32'b00000000000000010101001011011111; // input=-0.88037109375, output=2.64744038691
			11'd1926: out = 32'b00000000000000010101001100100011; // input=-0.88134765625, output=2.64950335647
			11'd1927: out = 32'b00000000000000010101001101100111; // input=-0.88232421875, output=2.65157429567
			11'd1928: out = 32'b00000000000000010101001110101011; // input=-0.88330078125, output=2.65365330659
			11'd1929: out = 32'b00000000000000010101001111101111; // input=-0.88427734375, output=2.65574049343
			11'd1930: out = 32'b00000000000000010101010000110100; // input=-0.88525390625, output=2.65783596262
			11'd1931: out = 32'b00000000000000010101010001111001; // input=-0.88623046875, output=2.65993982287
			11'd1932: out = 32'b00000000000000010101010010111110; // input=-0.88720703125, output=2.66205218521
			11'd1933: out = 32'b00000000000000010101010100000100; // input=-0.88818359375, output=2.6641731631
			11'd1934: out = 32'b00000000000000010101010101001001; // input=-0.88916015625, output=2.66630287249
			11'd1935: out = 32'b00000000000000010101010110001111; // input=-0.89013671875, output=2.6684414319
			11'd1936: out = 32'b00000000000000010101010111010110; // input=-0.89111328125, output=2.67058896248
			11'd1937: out = 32'b00000000000000010101011000011101; // input=-0.89208984375, output=2.67274558811
			11'd1938: out = 32'b00000000000000010101011001100011; // input=-0.89306640625, output=2.67491143551
			11'd1939: out = 32'b00000000000000010101011010101011; // input=-0.89404296875, output=2.67708663428
			11'd1940: out = 32'b00000000000000010101011011110010; // input=-0.89501953125, output=2.67927131704
			11'd1941: out = 32'b00000000000000010101011100111010; // input=-0.89599609375, output=2.6814656195
			11'd1942: out = 32'b00000000000000010101011110000010; // input=-0.89697265625, output=2.68366968056
			11'd1943: out = 32'b00000000000000010101011111001011; // input=-0.89794921875, output=2.68588364245
			11'd1944: out = 32'b00000000000000010101100000010100; // input=-0.89892578125, output=2.6881076508
			11'd1945: out = 32'b00000000000000010101100001011101; // input=-0.89990234375, output=2.69034185478
			11'd1946: out = 32'b00000000000000010101100010100111; // input=-0.90087890625, output=2.69258640723
			11'd1947: out = 32'b00000000000000010101100011110001; // input=-0.90185546875, output=2.69484146476
			11'd1948: out = 32'b00000000000000010101100100111011; // input=-0.90283203125, output=2.69710718789
			11'd1949: out = 32'b00000000000000010101100110000101; // input=-0.90380859375, output=2.6993837412
			11'd1950: out = 32'b00000000000000010101100111010000; // input=-0.90478515625, output=2.70167129347
			11'd1951: out = 32'b00000000000000010101101000011100; // input=-0.90576171875, output=2.70397001782
			11'd1952: out = 32'b00000000000000010101101001100111; // input=-0.90673828125, output=2.70628009189
			11'd1953: out = 32'b00000000000000010101101010110011; // input=-0.90771484375, output=2.70860169798
			11'd1954: out = 32'b00000000000000010101101100000000; // input=-0.90869140625, output=2.71093502324
			11'd1955: out = 32'b00000000000000010101101101001101; // input=-0.90966796875, output=2.71328025987
			11'd1956: out = 32'b00000000000000010101101110011010; // input=-0.91064453125, output=2.71563760525
			11'd1957: out = 32'b00000000000000010101101111101000; // input=-0.91162109375, output=2.71800726222
			11'd1958: out = 32'b00000000000000010101110000110110; // input=-0.91259765625, output=2.72038943924
			11'd1959: out = 32'b00000000000000010101110010000100; // input=-0.91357421875, output=2.72278435059
			11'd1960: out = 32'b00000000000000010101110011010011; // input=-0.91455078125, output=2.72519221669
			11'd1961: out = 32'b00000000000000010101110100100010; // input=-0.91552734375, output=2.72761326425
			11'd1962: out = 32'b00000000000000010101110101110010; // input=-0.91650390625, output=2.73004772657
			11'd1963: out = 32'b00000000000000010101110111000010; // input=-0.91748046875, output=2.73249584383
			11'd1964: out = 32'b00000000000000010101111000010011; // input=-0.91845703125, output=2.73495786332
			11'd1965: out = 32'b00000000000000010101111001100100; // input=-0.91943359375, output=2.73743403981
			11'd1966: out = 32'b00000000000000010101111010110110; // input=-0.92041015625, output=2.73992463579
			11'd1967: out = 32'b00000000000000010101111100001000; // input=-0.92138671875, output=2.74242992187
			11'd1968: out = 32'b00000000000000010101111101011011; // input=-0.92236328125, output=2.74495017711
			11'd1969: out = 32'b00000000000000010101111110101110; // input=-0.92333984375, output=2.74748568938
			11'd1970: out = 32'b00000000000000010110000000000001; // input=-0.92431640625, output=2.75003675577
			11'd1971: out = 32'b00000000000000010110000001010101; // input=-0.92529296875, output=2.752603683
			11'd1972: out = 32'b00000000000000010110000010101010; // input=-0.92626953125, output=2.75518678789
			11'd1973: out = 32'b00000000000000010110000011111111; // input=-0.92724609375, output=2.75778639778
			11'd1974: out = 32'b00000000000000010110000101010101; // input=-0.92822265625, output=2.76040285107
			11'd1975: out = 32'b00000000000000010110000110101011; // input=-0.92919921875, output=2.76303649773
			11'd1976: out = 32'b00000000000000010110001000000010; // input=-0.93017578125, output=2.76568769986
			11'd1977: out = 32'b00000000000000010110001001011010; // input=-0.93115234375, output=2.76835683229
			11'd1978: out = 32'b00000000000000010110001010110010; // input=-0.93212890625, output=2.77104428323
			11'd1979: out = 32'b00000000000000010110001100001010; // input=-0.93310546875, output=2.77375045491
			11'd1980: out = 32'b00000000000000010110001101100100; // input=-0.93408203125, output=2.77647576435
			11'd1981: out = 32'b00000000000000010110001110111110; // input=-0.93505859375, output=2.77922064407
			11'd1982: out = 32'b00000000000000010110010000011000; // input=-0.93603515625, output=2.78198554298
			11'd1983: out = 32'b00000000000000010110010001110011; // input=-0.93701171875, output=2.7847709272
			11'd1984: out = 32'b00000000000000010110010011001111; // input=-0.93798828125, output=2.78757728101
			11'd1985: out = 32'b00000000000000010110010100101100; // input=-0.93896484375, output=2.79040510791
			11'd1986: out = 32'b00000000000000010110010110001001; // input=-0.93994140625, output=2.79325493161
			11'd1987: out = 32'b00000000000000010110010111100111; // input=-0.94091796875, output=2.79612729726
			11'd1988: out = 32'b00000000000000010110011001000110; // input=-0.94189453125, output=2.79902277268
			11'd1989: out = 32'b00000000000000010110011010100110; // input=-0.94287109375, output=2.80194194967
			11'd1990: out = 32'b00000000000000010110011100000110; // input=-0.94384765625, output=2.8048854455
			11'd1991: out = 32'b00000000000000010110011101101000; // input=-0.94482421875, output=2.80785390442
			11'd1992: out = 32'b00000000000000010110011111001010; // input=-0.94580078125, output=2.81084799938
			11'd1993: out = 32'b00000000000000010110100000101101; // input=-0.94677734375, output=2.81386843382
			11'd1994: out = 32'b00000000000000010110100010010001; // input=-0.94775390625, output=2.81691594366
			11'd1995: out = 32'b00000000000000010110100011110101; // input=-0.94873046875, output=2.81999129943
			11'd1996: out = 32'b00000000000000010110100101011011; // input=-0.94970703125, output=2.8230953086
			11'd1997: out = 32'b00000000000000010110100111000010; // input=-0.95068359375, output=2.82622881808
			11'd1998: out = 32'b00000000000000010110101000101010; // input=-0.95166015625, output=2.82939271698
			11'd1999: out = 32'b00000000000000010110101010010010; // input=-0.95263671875, output=2.83258793963
			11'd2000: out = 32'b00000000000000010110101011111100; // input=-0.95361328125, output=2.83581546885
			11'd2001: out = 32'b00000000000000010110101101100111; // input=-0.95458984375, output=2.83907633955
			11'd2002: out = 32'b00000000000000010110101111010011; // input=-0.95556640625, output=2.84237164265
			11'd2003: out = 32'b00000000000000010110110001000000; // input=-0.95654296875, output=2.84570252945
			11'd2004: out = 32'b00000000000000010110110010101110; // input=-0.95751953125, output=2.84907021641
			11'd2005: out = 32'b00000000000000010110110100011110; // input=-0.95849609375, output=2.85247599038
			11'd2006: out = 32'b00000000000000010110110110001111; // input=-0.95947265625, output=2.85592121451
			11'd2007: out = 32'b00000000000000010110111000000001; // input=-0.96044921875, output=2.85940733468
			11'd2008: out = 32'b00000000000000010110111001110101; // input=-0.96142578125, output=2.86293588669
			11'd2009: out = 32'b00000000000000010110111011101010; // input=-0.96240234375, output=2.86650850434
			11'd2010: out = 32'b00000000000000010110111101100000; // input=-0.96337890625, output=2.87012692836
			11'd2011: out = 32'b00000000000000010110111111011000; // input=-0.96435546875, output=2.87379301647
			11'd2012: out = 32'b00000000000000010111000001010010; // input=-0.96533203125, output=2.87750875471
			11'd2013: out = 32'b00000000000000010111000011001110; // input=-0.96630859375, output=2.88127627019
			11'd2014: out = 32'b00000000000000010111000101001011; // input=-0.96728515625, output=2.88509784549
			11'd2015: out = 32'b00000000000000010111000111001010; // input=-0.96826171875, output=2.88897593506
			11'd2016: out = 32'b00000000000000010111001001001011; // input=-0.96923828125, output=2.89291318391
			11'd2017: out = 32'b00000000000000010111001011001110; // input=-0.97021484375, output=2.89691244895
			11'd2018: out = 32'b00000000000000010111001101010011; // input=-0.97119140625, output=2.90097682353
			11'd2019: out = 32'b00000000000000010111001111011011; // input=-0.97216796875, output=2.90510966579
			11'd2020: out = 32'b00000000000000010111010001100100; // input=-0.97314453125, output=2.90931463147
			11'd2021: out = 32'b00000000000000010111010011110001; // input=-0.97412109375, output=2.91359571221
			11'd2022: out = 32'b00000000000000010111010110000000; // input=-0.97509765625, output=2.91795728034
			11'd2023: out = 32'b00000000000000010111011000010001; // input=-0.97607421875, output=2.92240414177
			11'd2024: out = 32'b00000000000000010111011010100110; // input=-0.97705078125, output=2.92694159862
			11'd2025: out = 32'b00000000000000010111011100111110; // input=-0.97802734375, output=2.93157552401
			11'd2026: out = 32'b00000000000000010111011111011001; // input=-0.97900390625, output=2.93631245203
			11'd2027: out = 32'b00000000000000010111100001111000; // input=-0.97998046875, output=2.94115968675
			11'd2028: out = 32'b00000000000000010111100100011011; // input=-0.98095703125, output=2.94612543553
			11'd2029: out = 32'b00000000000000010111100111000010; // input=-0.98193359375, output=2.95121897351
			11'd2030: out = 32'b00000000000000010111101001101101; // input=-0.98291015625, output=2.95645084881
			11'd2031: out = 32'b00000000000000010111101100011101; // input=-0.98388671875, output=2.9618331413
			11'd2032: out = 32'b00000000000000010111101111010011; // input=-0.98486328125, output=2.96737979326
			11'd2033: out = 32'b00000000000000010111110010001111; // input=-0.98583984375, output=2.97310703786
			11'd2034: out = 32'b00000000000000010111110101010001; // input=-0.98681640625, output=2.97903396338
			11'd2035: out = 32'b00000000000000010111111000011010; // input=-0.98779296875, output=2.98518326972
			11'd2036: out = 32'b00000000000000010111111011101100; // input=-0.98876953125, output=2.99158230393
			11'd2037: out = 32'b00000000000000010111111111000111; // input=-0.98974609375, output=2.99826451197
			11'd2038: out = 32'b00000000000000011000000010101101; // input=-0.99072265625, output=3.00527153127
			11'd2039: out = 32'b00000000000000011000000110011111; // input=-0.99169921875, output=3.01265630832
			11'd2040: out = 32'b00000000000000011000001010011111; // input=-0.99267578125, output=3.02048793072
			11'd2041: out = 32'b00000000000000011000001110110010; // input=-0.99365234375, output=3.0288594899
			11'd2042: out = 32'b00000000000000011000010011011010; // input=-0.99462890625, output=3.03790168237
			11'd2043: out = 32'b00000000000000011000011000011111; // input=-0.99560546875, output=3.04780828732
			11'd2044: out = 32'b00000000000000011000011110001010; // input=-0.99658203125, output=3.05888935726
			11'd2045: out = 32'b00000000000000011000100100101110; // input=-0.99755859375, output=3.07170130494
			11'd2046: out = 32'b00000000000000011000101100110010; // input=-0.99853515625, output=3.08745945643
			11'd2047: out = 32'b00000000000000011000111000100000; // input=-0.99951171875, output=3.11034138188
		endcase
	end
	converter_arc U0 (a, index);

endmodule
