// Developed by: 	Amir Yazdanbakhsh
// Email: 			a.yazdanbakhsh@gatech.edu

`timescale 1ns/1ps
module log_lut(d_in, d_out);
	input		[31:0] d_in;
	output	reg	[31:0] d_out;

	wire	[10:0] addr;

	always @(addr)
		begin:lut_rom
			case(addr)
				11'd0: d_out <= 32'b00000000000000000000000000000000; // d_in = 1.000000, d_out = 0.000000
				11'd1: d_out <= 32'b00000000000000000000000010000000; // d_in = 1.001953, d_out = 0.001951
				11'd2: d_out <= 32'b00000000000000000000000100000000; // d_in = 1.003906, d_out = 0.003899
				11'd3: d_out <= 32'b00000000000000000000000101111111; // d_in = 1.005859, d_out = 0.005842
				11'd4: d_out <= 32'b00000000000000000000000111111110; // d_in = 1.007812, d_out = 0.007782
				11'd5: d_out <= 32'b00000000000000000000001001111101; // d_in = 1.009766, d_out = 0.009718
				11'd6: d_out <= 32'b00000000000000000000001011111100; // d_in = 1.011719, d_out = 0.011651
				11'd7: d_out <= 32'b00000000000000000000001101111010; // d_in = 1.013672, d_out = 0.013579
				11'd8: d_out <= 32'b00000000000000000000001111111000; // d_in = 1.015625, d_out = 0.015504
				11'd9: d_out <= 32'b00000000000000000000010001110110; // d_in = 1.017578, d_out = 0.017425
				11'd10: d_out <= 32'b00000000000000000000010011110100; // d_in = 1.019531, d_out = 0.019343
				11'd11: d_out <= 32'b00000000000000000000010101110001; // d_in = 1.021484, d_out = 0.021257
				11'd12: d_out <= 32'b00000000000000000000010111101110; // d_in = 1.023438, d_out = 0.023167
				11'd13: d_out <= 32'b00000000000000000000011001101011; // d_in = 1.025391, d_out = 0.025074
				11'd14: d_out <= 32'b00000000000000000000011011101000; // d_in = 1.027344, d_out = 0.026977
				11'd15: d_out <= 32'b00000000000000000000011101100100; // d_in = 1.029297, d_out = 0.028876
				11'd16: d_out <= 32'b00000000000000000000011111100001; // d_in = 1.031250, d_out = 0.030772
				11'd17: d_out <= 32'b00000000000000000000100001011101; // d_in = 1.033203, d_out = 0.032664
				11'd18: d_out <= 32'b00000000000000000000100011011000; // d_in = 1.035156, d_out = 0.034552
				11'd19: d_out <= 32'b00000000000000000000100101010100; // d_in = 1.037109, d_out = 0.036437
				11'd20: d_out <= 32'b00000000000000000000100111001111; // d_in = 1.039062, d_out = 0.038319
				11'd21: d_out <= 32'b00000000000000000000101001001010; // d_in = 1.041016, d_out = 0.040197
				11'd22: d_out <= 32'b00000000000000000000101011000101; // d_in = 1.042969, d_out = 0.042071
				11'd23: d_out <= 32'b00000000000000000000101101000000; // d_in = 1.044922, d_out = 0.043942
				11'd24: d_out <= 32'b00000000000000000000101110111010; // d_in = 1.046875, d_out = 0.045810
				11'd25: d_out <= 32'b00000000000000000000110000110100; // d_in = 1.048828, d_out = 0.047673
				11'd26: d_out <= 32'b00000000000000000000110010101110; // d_in = 1.050781, d_out = 0.049534
				11'd27: d_out <= 32'b00000000000000000000110100101000; // d_in = 1.052734, d_out = 0.051391
				11'd28: d_out <= 32'b00000000000000000000110110100001; // d_in = 1.054688, d_out = 0.053245
				11'd29: d_out <= 32'b00000000000000000000111000011011; // d_in = 1.056641, d_out = 0.055095
				11'd30: d_out <= 32'b00000000000000000000111010010100; // d_in = 1.058594, d_out = 0.056941
				11'd31: d_out <= 32'b00000000000000000000111100001101; // d_in = 1.060547, d_out = 0.058785
				11'd32: d_out <= 32'b00000000000000000000111110000101; // d_in = 1.062500, d_out = 0.060625
				11'd33: d_out <= 32'b00000000000000000000111111111101; // d_in = 1.064453, d_out = 0.062461
				11'd34: d_out <= 32'b00000000000000000001000001110110; // d_in = 1.066406, d_out = 0.064294
				11'd35: d_out <= 32'b00000000000000000001000011101110; // d_in = 1.068359, d_out = 0.066124
				11'd36: d_out <= 32'b00000000000000000001000101100101; // d_in = 1.070312, d_out = 0.067951
				11'd37: d_out <= 32'b00000000000000000001000111011101; // d_in = 1.072266, d_out = 0.069774
				11'd38: d_out <= 32'b00000000000000000001001001010100; // d_in = 1.074219, d_out = 0.071594
				11'd39: d_out <= 32'b00000000000000000001001011001011; // d_in = 1.076172, d_out = 0.073410
				11'd40: d_out <= 32'b00000000000000000001001101000010; // d_in = 1.078125, d_out = 0.075223
				11'd41: d_out <= 32'b00000000000000000001001110111000; // d_in = 1.080078, d_out = 0.077033
				11'd42: d_out <= 32'b00000000000000000001010000101111; // d_in = 1.082031, d_out = 0.078840
				11'd43: d_out <= 32'b00000000000000000001010010100101; // d_in = 1.083984, d_out = 0.080643
				11'd44: d_out <= 32'b00000000000000000001010100011011; // d_in = 1.085938, d_out = 0.082444
				11'd45: d_out <= 32'b00000000000000000001010110010001; // d_in = 1.087891, d_out = 0.084241
				11'd46: d_out <= 32'b00000000000000000001011000000110; // d_in = 1.089844, d_out = 0.086034
				11'd47: d_out <= 32'b00000000000000000001011001111100; // d_in = 1.091797, d_out = 0.087825
				11'd48: d_out <= 32'b00000000000000000001011011110001; // d_in = 1.093750, d_out = 0.089612
				11'd49: d_out <= 32'b00000000000000000001011101100110; // d_in = 1.095703, d_out = 0.091396
				11'd50: d_out <= 32'b00000000000000000001011111011010; // d_in = 1.097656, d_out = 0.093177
				11'd51: d_out <= 32'b00000000000000000001100001001111; // d_in = 1.099609, d_out = 0.094955
				11'd52: d_out <= 32'b00000000000000000001100011000011; // d_in = 1.101562, d_out = 0.096730
				11'd53: d_out <= 32'b00000000000000000001100100110111; // d_in = 1.103516, d_out = 0.098501
				11'd54: d_out <= 32'b00000000000000000001100110101011; // d_in = 1.105469, d_out = 0.100269
				11'd55: d_out <= 32'b00000000000000000001101000011111; // d_in = 1.107422, d_out = 0.102035
				11'd56: d_out <= 32'b00000000000000000001101010010010; // d_in = 1.109375, d_out = 0.103797
				11'd57: d_out <= 32'b00000000000000000001101100000110; // d_in = 1.111328, d_out = 0.105556
				11'd58: d_out <= 32'b00000000000000000001101101111001; // d_in = 1.113281, d_out = 0.107312
				11'd59: d_out <= 32'b00000000000000000001101111101100; // d_in = 1.115234, d_out = 0.109065
				11'd60: d_out <= 32'b00000000000000000001110001011110; // d_in = 1.117188, d_out = 0.110814
				11'd61: d_out <= 32'b00000000000000000001110011010001; // d_in = 1.119141, d_out = 0.112561
				11'd62: d_out <= 32'b00000000000000000001110101000011; // d_in = 1.121094, d_out = 0.114305
				11'd63: d_out <= 32'b00000000000000000001110110110101; // d_in = 1.123047, d_out = 0.116045
				11'd64: d_out <= 32'b00000000000000000001111000100111; // d_in = 1.125000, d_out = 0.117783
				11'd65: d_out <= 32'b00000000000000000001111010011001; // d_in = 1.126953, d_out = 0.119518
				11'd66: d_out <= 32'b00000000000000000001111100001010; // d_in = 1.128906, d_out = 0.121249
				11'd67: d_out <= 32'b00000000000000000001111101111011; // d_in = 1.130859, d_out = 0.122978
				11'd68: d_out <= 32'b00000000000000000001111111101101; // d_in = 1.132812, d_out = 0.124703
				11'd69: d_out <= 32'b00000000000000000010000001011101; // d_in = 1.134766, d_out = 0.126426
				11'd70: d_out <= 32'b00000000000000000010000011001110; // d_in = 1.136719, d_out = 0.128146
				11'd71: d_out <= 32'b00000000000000000010000100111111; // d_in = 1.138672, d_out = 0.129863
				11'd72: d_out <= 32'b00000000000000000010000110101111; // d_in = 1.140625, d_out = 0.131576
				11'd73: d_out <= 32'b00000000000000000010001000011111; // d_in = 1.142578, d_out = 0.133287
				11'd74: d_out <= 32'b00000000000000000010001010001111; // d_in = 1.144531, d_out = 0.134995
				11'd75: d_out <= 32'b00000000000000000010001011111111; // d_in = 1.146484, d_out = 0.136700
				11'd76: d_out <= 32'b00000000000000000010001101101110; // d_in = 1.148438, d_out = 0.138402
				11'd77: d_out <= 32'b00000000000000000010001111011110; // d_in = 1.150391, d_out = 0.140102
				11'd78: d_out <= 32'b00000000000000000010010001001101; // d_in = 1.152344, d_out = 0.141798
				11'd79: d_out <= 32'b00000000000000000010010010111100; // d_in = 1.154297, d_out = 0.143491
				11'd80: d_out <= 32'b00000000000000000010010100101011; // d_in = 1.156250, d_out = 0.145182
				11'd81: d_out <= 32'b00000000000000000010010110011001; // d_in = 1.158203, d_out = 0.146870
				11'd82: d_out <= 32'b00000000000000000010011000001000; // d_in = 1.160156, d_out = 0.148555
				11'd83: d_out <= 32'b00000000000000000010011001110110; // d_in = 1.162109, d_out = 0.150237
				11'd84: d_out <= 32'b00000000000000000010011011100100; // d_in = 1.164062, d_out = 0.151916
				11'd85: d_out <= 32'b00000000000000000010011101010010; // d_in = 1.166016, d_out = 0.153592
				11'd86: d_out <= 32'b00000000000000000010011111000000; // d_in = 1.167969, d_out = 0.155266
				11'd87: d_out <= 32'b00000000000000000010100000101101; // d_in = 1.169922, d_out = 0.156937
				11'd88: d_out <= 32'b00000000000000000010100010011010; // d_in = 1.171875, d_out = 0.158605
				11'd89: d_out <= 32'b00000000000000000010100100000111; // d_in = 1.173828, d_out = 0.160270
				11'd90: d_out <= 32'b00000000000000000010100101110100; // d_in = 1.175781, d_out = 0.161933
				11'd91: d_out <= 32'b00000000000000000010100111100001; // d_in = 1.177734, d_out = 0.163593
				11'd92: d_out <= 32'b00000000000000000010101001001110; // d_in = 1.179688, d_out = 0.165250
				11'd93: d_out <= 32'b00000000000000000010101010111010; // d_in = 1.181641, d_out = 0.166904
				11'd94: d_out <= 32'b00000000000000000010101100100110; // d_in = 1.183594, d_out = 0.168555
				11'd95: d_out <= 32'b00000000000000000010101110010011; // d_in = 1.185547, d_out = 0.170204
				11'd96: d_out <= 32'b00000000000000000010101111111110; // d_in = 1.187500, d_out = 0.171850
				11'd97: d_out <= 32'b00000000000000000010110001101010; // d_in = 1.189453, d_out = 0.173494
				11'd98: d_out <= 32'b00000000000000000010110011010110; // d_in = 1.191406, d_out = 0.175134
				11'd99: d_out <= 32'b00000000000000000010110101000001; // d_in = 1.193359, d_out = 0.176772
				11'd100: d_out <= 32'b00000000000000000010110110101100; // d_in = 1.195312, d_out = 0.178408
				11'd101: d_out <= 32'b00000000000000000010111000010111; // d_in = 1.197266, d_out = 0.180040
				11'd102: d_out <= 32'b00000000000000000010111010000010; // d_in = 1.199219, d_out = 0.181670
				11'd103: d_out <= 32'b00000000000000000010111011101101; // d_in = 1.201172, d_out = 0.183298
				11'd104: d_out <= 32'b00000000000000000010111101010111; // d_in = 1.203125, d_out = 0.184922
				11'd105: d_out <= 32'b00000000000000000010111111000001; // d_in = 1.205078, d_out = 0.186544
				11'd106: d_out <= 32'b00000000000000000011000000101100; // d_in = 1.207031, d_out = 0.188164
				11'd107: d_out <= 32'b00000000000000000011000010010101; // d_in = 1.208984, d_out = 0.189781
				11'd108: d_out <= 32'b00000000000000000011000011111111; // d_in = 1.210938, d_out = 0.191395
				11'd109: d_out <= 32'b00000000000000000011000101101001; // d_in = 1.212891, d_out = 0.193006
				11'd110: d_out <= 32'b00000000000000000011000111010010; // d_in = 1.214844, d_out = 0.194615
				11'd111: d_out <= 32'b00000000000000000011001000111100; // d_in = 1.216797, d_out = 0.196222
				11'd112: d_out <= 32'b00000000000000000011001010100101; // d_in = 1.218750, d_out = 0.197826
				11'd113: d_out <= 32'b00000000000000000011001100001110; // d_in = 1.220703, d_out = 0.199427
				11'd114: d_out <= 32'b00000000000000000011001101110110; // d_in = 1.222656, d_out = 0.201026
				11'd115: d_out <= 32'b00000000000000000011001111011111; // d_in = 1.224609, d_out = 0.202622
				11'd116: d_out <= 32'b00000000000000000011010001000111; // d_in = 1.226562, d_out = 0.204216
				11'd117: d_out <= 32'b00000000000000000011010010110000; // d_in = 1.228516, d_out = 0.205807
				11'd118: d_out <= 32'b00000000000000000011010100011000; // d_in = 1.230469, d_out = 0.207395
				11'd119: d_out <= 32'b00000000000000000011010110000000; // d_in = 1.232422, d_out = 0.208981
				11'd120: d_out <= 32'b00000000000000000011010111101000; // d_in = 1.234375, d_out = 0.210565
				11'd121: d_out <= 32'b00000000000000000011011001001111; // d_in = 1.236328, d_out = 0.212146
				11'd122: d_out <= 32'b00000000000000000011011010110111; // d_in = 1.238281, d_out = 0.213724
				11'd123: d_out <= 32'b00000000000000000011011100011110; // d_in = 1.240234, d_out = 0.215300
				11'd124: d_out <= 32'b00000000000000000011011110000101; // d_in = 1.242188, d_out = 0.216874
				11'd125: d_out <= 32'b00000000000000000011011111101100; // d_in = 1.244141, d_out = 0.218445
				11'd126: d_out <= 32'b00000000000000000011100001010011; // d_in = 1.246094, d_out = 0.220014
				11'd127: d_out <= 32'b00000000000000000011100010111001; // d_in = 1.248047, d_out = 0.221580
				11'd128: d_out <= 32'b00000000000000000011100100100000; // d_in = 1.250000, d_out = 0.223144
				11'd129: d_out <= 32'b00000000000000000011100110000110; // d_in = 1.251953, d_out = 0.224705
				11'd130: d_out <= 32'b00000000000000000011100111101100; // d_in = 1.253906, d_out = 0.226264
				11'd131: d_out <= 32'b00000000000000000011101001010010; // d_in = 1.255859, d_out = 0.227820
				11'd132: d_out <= 32'b00000000000000000011101010111000; // d_in = 1.257812, d_out = 0.229374
				11'd133: d_out <= 32'b00000000000000000011101100011110; // d_in = 1.259766, d_out = 0.230926
				11'd134: d_out <= 32'b00000000000000000011101110000011; // d_in = 1.261719, d_out = 0.232475
				11'd135: d_out <= 32'b00000000000000000011101111101001; // d_in = 1.263672, d_out = 0.234022
				11'd136: d_out <= 32'b00000000000000000011110001001110; // d_in = 1.265625, d_out = 0.235566
				11'd137: d_out <= 32'b00000000000000000011110010110011; // d_in = 1.267578, d_out = 0.237108
				11'd138: d_out <= 32'b00000000000000000011110100011000; // d_in = 1.269531, d_out = 0.238648
				11'd139: d_out <= 32'b00000000000000000011110101111101; // d_in = 1.271484, d_out = 0.240185
				11'd140: d_out <= 32'b00000000000000000011110111100001; // d_in = 1.273438, d_out = 0.241720
				11'd141: d_out <= 32'b00000000000000000011111001000110; // d_in = 1.275391, d_out = 0.243253
				11'd142: d_out <= 32'b00000000000000000011111010101010; // d_in = 1.277344, d_out = 0.244783
				11'd143: d_out <= 32'b00000000000000000011111100001110; // d_in = 1.279297, d_out = 0.246311
				11'd144: d_out <= 32'b00000000000000000011111101110010; // d_in = 1.281250, d_out = 0.247836
				11'd145: d_out <= 32'b00000000000000000011111111010110; // d_in = 1.283203, d_out = 0.249359
				11'd146: d_out <= 32'b00000000000000000100000000111010; // d_in = 1.285156, d_out = 0.250880
				11'd147: d_out <= 32'b00000000000000000100000010011101; // d_in = 1.287109, d_out = 0.252399
				11'd148: d_out <= 32'b00000000000000000100000100000001; // d_in = 1.289062, d_out = 0.253915
				11'd149: d_out <= 32'b00000000000000000100000101100100; // d_in = 1.291016, d_out = 0.255429
				11'd150: d_out <= 32'b00000000000000000100000111000111; // d_in = 1.292969, d_out = 0.256941
				11'd151: d_out <= 32'b00000000000000000100001000101010; // d_in = 1.294922, d_out = 0.258450
				11'd152: d_out <= 32'b00000000000000000100001010001101; // d_in = 1.296875, d_out = 0.259958
				11'd153: d_out <= 32'b00000000000000000100001011101111; // d_in = 1.298828, d_out = 0.261462
				11'd154: d_out <= 32'b00000000000000000100001101010010; // d_in = 1.300781, d_out = 0.262965
				11'd155: d_out <= 32'b00000000000000000100001110110100; // d_in = 1.302734, d_out = 0.264465
				11'd156: d_out <= 32'b00000000000000000100010000010110; // d_in = 1.304688, d_out = 0.265964
				11'd157: d_out <= 32'b00000000000000000100010001111000; // d_in = 1.306641, d_out = 0.267459
				11'd158: d_out <= 32'b00000000000000000100010011011010; // d_in = 1.308594, d_out = 0.268953
				11'd159: d_out <= 32'b00000000000000000100010100111100; // d_in = 1.310547, d_out = 0.270445
				11'd160: d_out <= 32'b00000000000000000100010110011101; // d_in = 1.312500, d_out = 0.271934
				11'd161: d_out <= 32'b00000000000000000100010111111111; // d_in = 1.314453, d_out = 0.273421
				11'd162: d_out <= 32'b00000000000000000100011001100000; // d_in = 1.316406, d_out = 0.274905
				11'd163: d_out <= 32'b00000000000000000100011011000001; // d_in = 1.318359, d_out = 0.276388
				11'd164: d_out <= 32'b00000000000000000100011100100010; // d_in = 1.320312, d_out = 0.277868
				11'd165: d_out <= 32'b00000000000000000100011110000011; // d_in = 1.322266, d_out = 0.279347
				11'd166: d_out <= 32'b00000000000000000100011111100100; // d_in = 1.324219, d_out = 0.280823
				11'd167: d_out <= 32'b00000000000000000100100001000101; // d_in = 1.326172, d_out = 0.282297
				11'd168: d_out <= 32'b00000000000000000100100010100101; // d_in = 1.328125, d_out = 0.283768
				11'd169: d_out <= 32'b00000000000000000100100100000101; // d_in = 1.330078, d_out = 0.285238
				11'd170: d_out <= 32'b00000000000000000100100101100110; // d_in = 1.332031, d_out = 0.286705
				11'd171: d_out <= 32'b00000000000000000100100111000110; // d_in = 1.333984, d_out = 0.288170
				11'd172: d_out <= 32'b00000000000000000100101000100101; // d_in = 1.335938, d_out = 0.289633
				11'd173: d_out <= 32'b00000000000000000100101010000101; // d_in = 1.337891, d_out = 0.291094
				11'd174: d_out <= 32'b00000000000000000100101011100101; // d_in = 1.339844, d_out = 0.292553
				11'd175: d_out <= 32'b00000000000000000100101101000100; // d_in = 1.341797, d_out = 0.294010
				11'd176: d_out <= 32'b00000000000000000100101110100100; // d_in = 1.343750, d_out = 0.295464
				11'd177: d_out <= 32'b00000000000000000100110000000011; // d_in = 1.345703, d_out = 0.296917
				11'd178: d_out <= 32'b00000000000000000100110001100010; // d_in = 1.347656, d_out = 0.298367
				11'd179: d_out <= 32'b00000000000000000100110011000001; // d_in = 1.349609, d_out = 0.299815
				11'd180: d_out <= 32'b00000000000000000100110100011111; // d_in = 1.351562, d_out = 0.301261
				11'd181: d_out <= 32'b00000000000000000100110101111110; // d_in = 1.353516, d_out = 0.302705
				11'd182: d_out <= 32'b00000000000000000100110111011101; // d_in = 1.355469, d_out = 0.304147
				11'd183: d_out <= 32'b00000000000000000100111000111011; // d_in = 1.357422, d_out = 0.305587
				11'd184: d_out <= 32'b00000000000000000100111010011001; // d_in = 1.359375, d_out = 0.307025
				11'd185: d_out <= 32'b00000000000000000100111011110111; // d_in = 1.361328, d_out = 0.308461
				11'd186: d_out <= 32'b00000000000000000100111101010101; // d_in = 1.363281, d_out = 0.309894
				11'd187: d_out <= 32'b00000000000000000100111110110011; // d_in = 1.365234, d_out = 0.311326
				11'd188: d_out <= 32'b00000000000000000101000000010001; // d_in = 1.367188, d_out = 0.312756
				11'd189: d_out <= 32'b00000000000000000101000001101110; // d_in = 1.369141, d_out = 0.314183
				11'd190: d_out <= 32'b00000000000000000101000011001100; // d_in = 1.371094, d_out = 0.315609
				11'd191: d_out <= 32'b00000000000000000101000100101001; // d_in = 1.373047, d_out = 0.317032
				11'd192: d_out <= 32'b00000000000000000101000110000110; // d_in = 1.375000, d_out = 0.318454
				11'd193: d_out <= 32'b00000000000000000101000111100011; // d_in = 1.376953, d_out = 0.319873
				11'd194: d_out <= 32'b00000000000000000101001001000000; // d_in = 1.378906, d_out = 0.321291
				11'd195: d_out <= 32'b00000000000000000101001010011101; // d_in = 1.380859, d_out = 0.322706
				11'd196: d_out <= 32'b00000000000000000101001011111001; // d_in = 1.382812, d_out = 0.324119
				11'd197: d_out <= 32'b00000000000000000101001101010110; // d_in = 1.384766, d_out = 0.325531
				11'd198: d_out <= 32'b00000000000000000101001110110010; // d_in = 1.386719, d_out = 0.326940
				11'd199: d_out <= 32'b00000000000000000101010000001111; // d_in = 1.388672, d_out = 0.328348
				11'd200: d_out <= 32'b00000000000000000101010001101011; // d_in = 1.390625, d_out = 0.329753
				11'd201: d_out <= 32'b00000000000000000101010011000111; // d_in = 1.392578, d_out = 0.331157
				11'd202: d_out <= 32'b00000000000000000101010100100011; // d_in = 1.394531, d_out = 0.332558
				11'd203: d_out <= 32'b00000000000000000101010101111110; // d_in = 1.396484, d_out = 0.333958
				11'd204: d_out <= 32'b00000000000000000101010111011010; // d_in = 1.398438, d_out = 0.335356
				11'd205: d_out <= 32'b00000000000000000101011000110101; // d_in = 1.400391, d_out = 0.336751
				11'd206: d_out <= 32'b00000000000000000101011010010001; // d_in = 1.402344, d_out = 0.338145
				11'd207: d_out <= 32'b00000000000000000101011011101100; // d_in = 1.404297, d_out = 0.339537
				11'd208: d_out <= 32'b00000000000000000101011101000111; // d_in = 1.406250, d_out = 0.340927
				11'd209: d_out <= 32'b00000000000000000101011110100010; // d_in = 1.408203, d_out = 0.342315
				11'd210: d_out <= 32'b00000000000000000101011111111101; // d_in = 1.410156, d_out = 0.343701
				11'd211: d_out <= 32'b00000000000000000101100001010111; // d_in = 1.412109, d_out = 0.345085
				11'd212: d_out <= 32'b00000000000000000101100010110010; // d_in = 1.414062, d_out = 0.346467
				11'd213: d_out <= 32'b00000000000000000101100100001101; // d_in = 1.416016, d_out = 0.347847
				11'd214: d_out <= 32'b00000000000000000101100101100111; // d_in = 1.417969, d_out = 0.349225
				11'd215: d_out <= 32'b00000000000000000101100111000001; // d_in = 1.419922, d_out = 0.350602
				11'd216: d_out <= 32'b00000000000000000101101000011011; // d_in = 1.421875, d_out = 0.351976
				11'd217: d_out <= 32'b00000000000000000101101001110101; // d_in = 1.423828, d_out = 0.353349
				11'd218: d_out <= 32'b00000000000000000101101011001111; // d_in = 1.425781, d_out = 0.354720
				11'd219: d_out <= 32'b00000000000000000101101100101001; // d_in = 1.427734, d_out = 0.356089
				11'd220: d_out <= 32'b00000000000000000101101110000010; // d_in = 1.429688, d_out = 0.357456
				11'd221: d_out <= 32'b00000000000000000101101111011100; // d_in = 1.431641, d_out = 0.358821
				11'd222: d_out <= 32'b00000000000000000101110000110101; // d_in = 1.433594, d_out = 0.360184
				11'd223: d_out <= 32'b00000000000000000101110010001110; // d_in = 1.435547, d_out = 0.361546
				11'd224: d_out <= 32'b00000000000000000101110011100111; // d_in = 1.437500, d_out = 0.362905
				11'd225: d_out <= 32'b00000000000000000101110101000000; // d_in = 1.439453, d_out = 0.364263
				11'd226: d_out <= 32'b00000000000000000101110110011001; // d_in = 1.441406, d_out = 0.365619
				11'd227: d_out <= 32'b00000000000000000101110111110010; // d_in = 1.443359, d_out = 0.366973
				11'd228: d_out <= 32'b00000000000000000101111001001011; // d_in = 1.445312, d_out = 0.368326
				11'd229: d_out <= 32'b00000000000000000101111010100011; // d_in = 1.447266, d_out = 0.369676
				11'd230: d_out <= 32'b00000000000000000101111011111011; // d_in = 1.449219, d_out = 0.371025
				11'd231: d_out <= 32'b00000000000000000101111101010100; // d_in = 1.451172, d_out = 0.372371
				11'd232: d_out <= 32'b00000000000000000101111110101100; // d_in = 1.453125, d_out = 0.373716
				11'd233: d_out <= 32'b00000000000000000110000000000100; // d_in = 1.455078, d_out = 0.375060
				11'd234: d_out <= 32'b00000000000000000110000001011100; // d_in = 1.457031, d_out = 0.376401
				11'd235: d_out <= 32'b00000000000000000110000010110100; // d_in = 1.458984, d_out = 0.377741
				11'd236: d_out <= 32'b00000000000000000110000100001011; // d_in = 1.460938, d_out = 0.379078
				11'd237: d_out <= 32'b00000000000000000110000101100011; // d_in = 1.462891, d_out = 0.380414
				11'd238: d_out <= 32'b00000000000000000110000110111010; // d_in = 1.464844, d_out = 0.381749
				11'd239: d_out <= 32'b00000000000000000110001000010010; // d_in = 1.466797, d_out = 0.383081
				11'd240: d_out <= 32'b00000000000000000110001001101001; // d_in = 1.468750, d_out = 0.384412
				11'd241: d_out <= 32'b00000000000000000110001011000000; // d_in = 1.470703, d_out = 0.385741
				11'd242: d_out <= 32'b00000000000000000110001100010111; // d_in = 1.472656, d_out = 0.387068
				11'd243: d_out <= 32'b00000000000000000110001101101110; // d_in = 1.474609, d_out = 0.388393
				11'd244: d_out <= 32'b00000000000000000110001111000100; // d_in = 1.476562, d_out = 0.389717
				11'd245: d_out <= 32'b00000000000000000110010000011011; // d_in = 1.478516, d_out = 0.391039
				11'd246: d_out <= 32'b00000000000000000110010001110010; // d_in = 1.480469, d_out = 0.392359
				11'd247: d_out <= 32'b00000000000000000110010011001000; // d_in = 1.482422, d_out = 0.393677
				11'd248: d_out <= 32'b00000000000000000110010100011110; // d_in = 1.484375, d_out = 0.394994
				11'd249: d_out <= 32'b00000000000000000110010101110100; // d_in = 1.486328, d_out = 0.396309
				11'd250: d_out <= 32'b00000000000000000110010111001011; // d_in = 1.488281, d_out = 0.397622
				11'd251: d_out <= 32'b00000000000000000110011000100000; // d_in = 1.490234, d_out = 0.398933
				11'd252: d_out <= 32'b00000000000000000110011001110110; // d_in = 1.492188, d_out = 0.400243
				11'd253: d_out <= 32'b00000000000000000110011011001100; // d_in = 1.494141, d_out = 0.401551
				11'd254: d_out <= 32'b00000000000000000110011100100010; // d_in = 1.496094, d_out = 0.402858
				11'd255: d_out <= 32'b00000000000000000110011101110111; // d_in = 1.498047, d_out = 0.404162
				11'd256: d_out <= 32'b00000000000000000110011111001101; // d_in = 1.500000, d_out = 0.405465
				11'd257: d_out <= 32'b00000000000000000110100000100010; // d_in = 1.501953, d_out = 0.406766
				11'd258: d_out <= 32'b00000000000000000110100001110111; // d_in = 1.503906, d_out = 0.408066
				11'd259: d_out <= 32'b00000000000000000110100011001100; // d_in = 1.505859, d_out = 0.409364
				11'd260: d_out <= 32'b00000000000000000110100100100001; // d_in = 1.507812, d_out = 0.410660
				11'd261: d_out <= 32'b00000000000000000110100101110110; // d_in = 1.509766, d_out = 0.411954
				11'd262: d_out <= 32'b00000000000000000110100111001011; // d_in = 1.511719, d_out = 0.413247
				11'd263: d_out <= 32'b00000000000000000110101000011111; // d_in = 1.513672, d_out = 0.414538
				11'd264: d_out <= 32'b00000000000000000110101001110100; // d_in = 1.515625, d_out = 0.415828
				11'd265: d_out <= 32'b00000000000000000110101011001000; // d_in = 1.517578, d_out = 0.417116
				11'd266: d_out <= 32'b00000000000000000110101100011100; // d_in = 1.519531, d_out = 0.418402
				11'd267: d_out <= 32'b00000000000000000110101101110001; // d_in = 1.521484, d_out = 0.419686
				11'd268: d_out <= 32'b00000000000000000110101111000101; // d_in = 1.523438, d_out = 0.420969
				11'd269: d_out <= 32'b00000000000000000110110000011001; // d_in = 1.525391, d_out = 0.422251
				11'd270: d_out <= 32'b00000000000000000110110001101100; // d_in = 1.527344, d_out = 0.423530
				11'd271: d_out <= 32'b00000000000000000110110011000000; // d_in = 1.529297, d_out = 0.424808
				11'd272: d_out <= 32'b00000000000000000110110100010100; // d_in = 1.531250, d_out = 0.426084
				11'd273: d_out <= 32'b00000000000000000110110101100111; // d_in = 1.533203, d_out = 0.427359
				11'd274: d_out <= 32'b00000000000000000110110110111011; // d_in = 1.535156, d_out = 0.428632
				11'd275: d_out <= 32'b00000000000000000110111000001110; // d_in = 1.537109, d_out = 0.429904
				11'd276: d_out <= 32'b00000000000000000110111001100001; // d_in = 1.539062, d_out = 0.431173
				11'd277: d_out <= 32'b00000000000000000110111010110100; // d_in = 1.541016, d_out = 0.432442
				11'd278: d_out <= 32'b00000000000000000110111100001000; // d_in = 1.542969, d_out = 0.433708
				11'd279: d_out <= 32'b00000000000000000110111101011010; // d_in = 1.544922, d_out = 0.434973
				11'd280: d_out <= 32'b00000000000000000110111110101101; // d_in = 1.546875, d_out = 0.436237
				11'd281: d_out <= 32'b00000000000000000111000000000000; // d_in = 1.548828, d_out = 0.437499
				11'd282: d_out <= 32'b00000000000000000111000001010010; // d_in = 1.550781, d_out = 0.438759
				11'd283: d_out <= 32'b00000000000000000111000010100101; // d_in = 1.552734, d_out = 0.440017
				11'd284: d_out <= 32'b00000000000000000111000011110111; // d_in = 1.554688, d_out = 0.441275
				11'd285: d_out <= 32'b00000000000000000111000101001010; // d_in = 1.556641, d_out = 0.442530
				11'd286: d_out <= 32'b00000000000000000111000110011100; // d_in = 1.558594, d_out = 0.443784
				11'd287: d_out <= 32'b00000000000000000111000111101110; // d_in = 1.560547, d_out = 0.445036
				11'd288: d_out <= 32'b00000000000000000111001001000000; // d_in = 1.562500, d_out = 0.446287
				11'd289: d_out <= 32'b00000000000000000111001010010010; // d_in = 1.564453, d_out = 0.447536
				11'd290: d_out <= 32'b00000000000000000111001011100100; // d_in = 1.566406, d_out = 0.448784
				11'd291: d_out <= 32'b00000000000000000111001100110101; // d_in = 1.568359, d_out = 0.450030
				11'd292: d_out <= 32'b00000000000000000111001110000111; // d_in = 1.570312, d_out = 0.451275
				11'd293: d_out <= 32'b00000000000000000111001111011000; // d_in = 1.572266, d_out = 0.452518
				11'd294: d_out <= 32'b00000000000000000111010000101010; // d_in = 1.574219, d_out = 0.453759
				11'd295: d_out <= 32'b00000000000000000111010001111011; // d_in = 1.576172, d_out = 0.454999
				11'd296: d_out <= 32'b00000000000000000111010011001100; // d_in = 1.578125, d_out = 0.456237
				11'd297: d_out <= 32'b00000000000000000111010100011101; // d_in = 1.580078, d_out = 0.457474
				11'd298: d_out <= 32'b00000000000000000111010101101110; // d_in = 1.582031, d_out = 0.458710
				11'd299: d_out <= 32'b00000000000000000111010110111111; // d_in = 1.583984, d_out = 0.459943
				11'd300: d_out <= 32'b00000000000000000111011000010000; // d_in = 1.585938, d_out = 0.461176
				11'd301: d_out <= 32'b00000000000000000111011001100000; // d_in = 1.587891, d_out = 0.462406
				11'd302: d_out <= 32'b00000000000000000111011010110001; // d_in = 1.589844, d_out = 0.463636
				11'd303: d_out <= 32'b00000000000000000111011100000001; // d_in = 1.591797, d_out = 0.464863
				11'd304: d_out <= 32'b00000000000000000111011101010010; // d_in = 1.593750, d_out = 0.466090
				11'd305: d_out <= 32'b00000000000000000111011110100010; // d_in = 1.595703, d_out = 0.467314
				11'd306: d_out <= 32'b00000000000000000111011111110010; // d_in = 1.597656, d_out = 0.468538
				11'd307: d_out <= 32'b00000000000000000111100001000010; // d_in = 1.599609, d_out = 0.469759
				11'd308: d_out <= 32'b00000000000000000111100010010010; // d_in = 1.601562, d_out = 0.470980
				11'd309: d_out <= 32'b00000000000000000111100011100010; // d_in = 1.603516, d_out = 0.472198
				11'd310: d_out <= 32'b00000000000000000111100100110010; // d_in = 1.605469, d_out = 0.473416
				11'd311: d_out <= 32'b00000000000000000111100110000001; // d_in = 1.607422, d_out = 0.474632
				11'd312: d_out <= 32'b00000000000000000111100111010001; // d_in = 1.609375, d_out = 0.475846
				11'd313: d_out <= 32'b00000000000000000111101000100001; // d_in = 1.611328, d_out = 0.477059
				11'd314: d_out <= 32'b00000000000000000111101001110000; // d_in = 1.613281, d_out = 0.478270
				11'd315: d_out <= 32'b00000000000000000111101010111111; // d_in = 1.615234, d_out = 0.479480
				11'd316: d_out <= 32'b00000000000000000111101100001110; // d_in = 1.617188, d_out = 0.480689
				11'd317: d_out <= 32'b00000000000000000111101101011110; // d_in = 1.619141, d_out = 0.481896
				11'd318: d_out <= 32'b00000000000000000111101110101101; // d_in = 1.621094, d_out = 0.483101
				11'd319: d_out <= 32'b00000000000000000111101111111011; // d_in = 1.623047, d_out = 0.484305
				11'd320: d_out <= 32'b00000000000000000111110001001010; // d_in = 1.625000, d_out = 0.485508
				11'd321: d_out <= 32'b00000000000000000111110010011001; // d_in = 1.626953, d_out = 0.486709
				11'd322: d_out <= 32'b00000000000000000111110011101000; // d_in = 1.628906, d_out = 0.487909
				11'd323: d_out <= 32'b00000000000000000111110100110110; // d_in = 1.630859, d_out = 0.489107
				11'd324: d_out <= 32'b00000000000000000111110110000101; // d_in = 1.632812, d_out = 0.490304
				11'd325: d_out <= 32'b00000000000000000111110111010011; // d_in = 1.634766, d_out = 0.491499
				11'd326: d_out <= 32'b00000000000000000111111000100001; // d_in = 1.636719, d_out = 0.492693
				11'd327: d_out <= 32'b00000000000000000111111001101111; // d_in = 1.638672, d_out = 0.493886
				11'd328: d_out <= 32'b00000000000000000111111010111101; // d_in = 1.640625, d_out = 0.495077
				11'd329: d_out <= 32'b00000000000000000111111100001011; // d_in = 1.642578, d_out = 0.496267
				11'd330: d_out <= 32'b00000000000000000111111101011001; // d_in = 1.644531, d_out = 0.497455
				11'd331: d_out <= 32'b00000000000000000111111110100111; // d_in = 1.646484, d_out = 0.498642
				11'd332: d_out <= 32'b00000000000000000111111111110101; // d_in = 1.648438, d_out = 0.499828
				11'd333: d_out <= 32'b00000000000000001000000001000010; // d_in = 1.650391, d_out = 0.501012
				11'd334: d_out <= 32'b00000000000000001000000010010000; // d_in = 1.652344, d_out = 0.502195
				11'd335: d_out <= 32'b00000000000000001000000011011101; // d_in = 1.654297, d_out = 0.503376
				11'd336: d_out <= 32'b00000000000000001000000100101011; // d_in = 1.656250, d_out = 0.504556
				11'd337: d_out <= 32'b00000000000000001000000101111000; // d_in = 1.658203, d_out = 0.505735
				11'd338: d_out <= 32'b00000000000000001000000111000101; // d_in = 1.660156, d_out = 0.506912
				11'd339: d_out <= 32'b00000000000000001000001000010010; // d_in = 1.662109, d_out = 0.508088
				11'd340: d_out <= 32'b00000000000000001000001001011111; // d_in = 1.664062, d_out = 0.509262
				11'd341: d_out <= 32'b00000000000000001000001010101100; // d_in = 1.666016, d_out = 0.510435
				11'd342: d_out <= 32'b00000000000000001000001011111001; // d_in = 1.667969, d_out = 0.511607
				11'd343: d_out <= 32'b00000000000000001000001101000101; // d_in = 1.669922, d_out = 0.512777
				11'd344: d_out <= 32'b00000000000000001000001110010010; // d_in = 1.671875, d_out = 0.513946
				11'd345: d_out <= 32'b00000000000000001000001111011110; // d_in = 1.673828, d_out = 0.515113
				11'd346: d_out <= 32'b00000000000000001000010000101011; // d_in = 1.675781, d_out = 0.516279
				11'd347: d_out <= 32'b00000000000000001000010001110111; // d_in = 1.677734, d_out = 0.517444
				11'd348: d_out <= 32'b00000000000000001000010011000011; // d_in = 1.679688, d_out = 0.518608
				11'd349: d_out <= 32'b00000000000000001000010100010000; // d_in = 1.681641, d_out = 0.519770
				11'd350: d_out <= 32'b00000000000000001000010101011100; // d_in = 1.683594, d_out = 0.520931
				11'd351: d_out <= 32'b00000000000000001000010110101000; // d_in = 1.685547, d_out = 0.522090
				11'd352: d_out <= 32'b00000000000000001000010111110100; // d_in = 1.687500, d_out = 0.523248
				11'd353: d_out <= 32'b00000000000000001000011000111111; // d_in = 1.689453, d_out = 0.524405
				11'd354: d_out <= 32'b00000000000000001000011010001011; // d_in = 1.691406, d_out = 0.525560
				11'd355: d_out <= 32'b00000000000000001000011011010111; // d_in = 1.693359, d_out = 0.526714
				11'd356: d_out <= 32'b00000000000000001000011100100010; // d_in = 1.695312, d_out = 0.527867
				11'd357: d_out <= 32'b00000000000000001000011101101110; // d_in = 1.697266, d_out = 0.529019
				11'd358: d_out <= 32'b00000000000000001000011110111001; // d_in = 1.699219, d_out = 0.530169
				11'd359: d_out <= 32'b00000000000000001000100000000100; // d_in = 1.701172, d_out = 0.531317
				11'd360: d_out <= 32'b00000000000000001000100001010000; // d_in = 1.703125, d_out = 0.532465
				11'd361: d_out <= 32'b00000000000000001000100010011011; // d_in = 1.705078, d_out = 0.533611
				11'd362: d_out <= 32'b00000000000000001000100011100110; // d_in = 1.707031, d_out = 0.534756
				11'd363: d_out <= 32'b00000000000000001000100100110001; // d_in = 1.708984, d_out = 0.535899
				11'd364: d_out <= 32'b00000000000000001000100101111100; // d_in = 1.710938, d_out = 0.537041
				11'd365: d_out <= 32'b00000000000000001000100111000110; // d_in = 1.712891, d_out = 0.538182
				11'd366: d_out <= 32'b00000000000000001000101000010001; // d_in = 1.714844, d_out = 0.539322
				11'd367: d_out <= 32'b00000000000000001000101001011100; // d_in = 1.716797, d_out = 0.540460
				11'd368: d_out <= 32'b00000000000000001000101010100110; // d_in = 1.718750, d_out = 0.541597
				11'd369: d_out <= 32'b00000000000000001000101011110001; // d_in = 1.720703, d_out = 0.542733
				11'd370: d_out <= 32'b00000000000000001000101100111011; // d_in = 1.722656, d_out = 0.543867
				11'd371: d_out <= 32'b00000000000000001000101110000101; // d_in = 1.724609, d_out = 0.545001
				11'd372: d_out <= 32'b00000000000000001000101111001111; // d_in = 1.726562, d_out = 0.546132
				11'd373: d_out <= 32'b00000000000000001000110000011001; // d_in = 1.728516, d_out = 0.547263
				11'd374: d_out <= 32'b00000000000000001000110001100011; // d_in = 1.730469, d_out = 0.548392
				11'd375: d_out <= 32'b00000000000000001000110010101101; // d_in = 1.732422, d_out = 0.549520
				11'd376: d_out <= 32'b00000000000000001000110011110111; // d_in = 1.734375, d_out = 0.550647
				11'd377: d_out <= 32'b00000000000000001000110101000001; // d_in = 1.736328, d_out = 0.551773
				11'd378: d_out <= 32'b00000000000000001000110110001011; // d_in = 1.738281, d_out = 0.552897
				11'd379: d_out <= 32'b00000000000000001000110111010100; // d_in = 1.740234, d_out = 0.554020
				11'd380: d_out <= 32'b00000000000000001000111000011110; // d_in = 1.742188, d_out = 0.555142
				11'd381: d_out <= 32'b00000000000000001000111001100111; // d_in = 1.744141, d_out = 0.556262
				11'd382: d_out <= 32'b00000000000000001000111010110001; // d_in = 1.746094, d_out = 0.557381
				11'd383: d_out <= 32'b00000000000000001000111011111010; // d_in = 1.748047, d_out = 0.558499
				11'd384: d_out <= 32'b00000000000000001000111101000011; // d_in = 1.750000, d_out = 0.559616
				11'd385: d_out <= 32'b00000000000000001000111110001100; // d_in = 1.751953, d_out = 0.560731
				11'd386: d_out <= 32'b00000000000000001000111111010101; // d_in = 1.753906, d_out = 0.561845
				11'd387: d_out <= 32'b00000000000000001001000000011110; // d_in = 1.755859, d_out = 0.562958
				11'd388: d_out <= 32'b00000000000000001001000001100111; // d_in = 1.757812, d_out = 0.564070
				11'd389: d_out <= 32'b00000000000000001001000010110000; // d_in = 1.759766, d_out = 0.565181
				11'd390: d_out <= 32'b00000000000000001001000011111000; // d_in = 1.761719, d_out = 0.566290
				11'd391: d_out <= 32'b00000000000000001001000101000001; // d_in = 1.763672, d_out = 0.567398
				11'd392: d_out <= 32'b00000000000000001001000110001010; // d_in = 1.765625, d_out = 0.568505
				11'd393: d_out <= 32'b00000000000000001001000111010010; // d_in = 1.767578, d_out = 0.569610
				11'd394: d_out <= 32'b00000000000000001001001000011010; // d_in = 1.769531, d_out = 0.570715
				11'd395: d_out <= 32'b00000000000000001001001001100011; // d_in = 1.771484, d_out = 0.571818
				11'd396: d_out <= 32'b00000000000000001001001010101011; // d_in = 1.773438, d_out = 0.572920
				11'd397: d_out <= 32'b00000000000000001001001011110011; // d_in = 1.775391, d_out = 0.574020
				11'd398: d_out <= 32'b00000000000000001001001100111011; // d_in = 1.777344, d_out = 0.575120
				11'd399: d_out <= 32'b00000000000000001001001110000011; // d_in = 1.779297, d_out = 0.576218
				11'd400: d_out <= 32'b00000000000000001001001111001011; // d_in = 1.781250, d_out = 0.577315
				11'd401: d_out <= 32'b00000000000000001001010000010011; // d_in = 1.783203, d_out = 0.578411
				11'd402: d_out <= 32'b00000000000000001001010001011011; // d_in = 1.785156, d_out = 0.579506
				11'd403: d_out <= 32'b00000000000000001001010010100010; // d_in = 1.787109, d_out = 0.580599
				11'd404: d_out <= 32'b00000000000000001001010011101010; // d_in = 1.789062, d_out = 0.581692
				11'd405: d_out <= 32'b00000000000000001001010100110001; // d_in = 1.791016, d_out = 0.582783
				11'd406: d_out <= 32'b00000000000000001001010101111001; // d_in = 1.792969, d_out = 0.583873
				11'd407: d_out <= 32'b00000000000000001001010111000000; // d_in = 1.794922, d_out = 0.584961
				11'd408: d_out <= 32'b00000000000000001001011000000111; // d_in = 1.796875, d_out = 0.586049
				11'd409: d_out <= 32'b00000000000000001001011001001111; // d_in = 1.798828, d_out = 0.587135
				11'd410: d_out <= 32'b00000000000000001001011010010110; // d_in = 1.800781, d_out = 0.588221
				11'd411: d_out <= 32'b00000000000000001001011011011101; // d_in = 1.802734, d_out = 0.589305
				11'd412: d_out <= 32'b00000000000000001001011100100100; // d_in = 1.804688, d_out = 0.590387
				11'd413: d_out <= 32'b00000000000000001001011101101011; // d_in = 1.806641, d_out = 0.591469
				11'd414: d_out <= 32'b00000000000000001001011110110001; // d_in = 1.808594, d_out = 0.592550
				11'd415: d_out <= 32'b00000000000000001001011111111000; // d_in = 1.810547, d_out = 0.593629
				11'd416: d_out <= 32'b00000000000000001001100000111111; // d_in = 1.812500, d_out = 0.594707
				11'd417: d_out <= 32'b00000000000000001001100010000101; // d_in = 1.814453, d_out = 0.595784
				11'd418: d_out <= 32'b00000000000000001001100011001100; // d_in = 1.816406, d_out = 0.596860
				11'd419: d_out <= 32'b00000000000000001001100100010010; // d_in = 1.818359, d_out = 0.597935
				11'd420: d_out <= 32'b00000000000000001001100101011001; // d_in = 1.820312, d_out = 0.599008
				11'd421: d_out <= 32'b00000000000000001001100110011111; // d_in = 1.822266, d_out = 0.600081
				11'd422: d_out <= 32'b00000000000000001001100111100101; // d_in = 1.824219, d_out = 0.601152
				11'd423: d_out <= 32'b00000000000000001001101000101011; // d_in = 1.826172, d_out = 0.602222
				11'd424: d_out <= 32'b00000000000000001001101001110001; // d_in = 1.828125, d_out = 0.603291
				11'd425: d_out <= 32'b00000000000000001001101010110111; // d_in = 1.830078, d_out = 0.604359
				11'd426: d_out <= 32'b00000000000000001001101011111101; // d_in = 1.832031, d_out = 0.605425
				11'd427: d_out <= 32'b00000000000000001001101101000011; // d_in = 1.833984, d_out = 0.606491
				11'd428: d_out <= 32'b00000000000000001001101110001001; // d_in = 1.835938, d_out = 0.607555
				11'd429: d_out <= 32'b00000000000000001001101111001110; // d_in = 1.837891, d_out = 0.608619
				11'd430: d_out <= 32'b00000000000000001001110000010100; // d_in = 1.839844, d_out = 0.609681
				11'd431: d_out <= 32'b00000000000000001001110001011010; // d_in = 1.841797, d_out = 0.610742
				11'd432: d_out <= 32'b00000000000000001001110010011111; // d_in = 1.843750, d_out = 0.611802
				11'd433: d_out <= 32'b00000000000000001001110011100100; // d_in = 1.845703, d_out = 0.612860
				11'd434: d_out <= 32'b00000000000000001001110100101010; // d_in = 1.847656, d_out = 0.613918
				11'd435: d_out <= 32'b00000000000000001001110101101111; // d_in = 1.849609, d_out = 0.614974
				11'd436: d_out <= 32'b00000000000000001001110110110100; // d_in = 1.851562, d_out = 0.616030
				11'd437: d_out <= 32'b00000000000000001001110111111001; // d_in = 1.853516, d_out = 0.617084
				11'd438: d_out <= 32'b00000000000000001001111000111110; // d_in = 1.855469, d_out = 0.618137
				11'd439: d_out <= 32'b00000000000000001001111010000011; // d_in = 1.857422, d_out = 0.619189
				11'd440: d_out <= 32'b00000000000000001001111011001000; // d_in = 1.859375, d_out = 0.620240
				11'd441: d_out <= 32'b00000000000000001001111100001101; // d_in = 1.861328, d_out = 0.621290
				11'd442: d_out <= 32'b00000000000000001001111101010010; // d_in = 1.863281, d_out = 0.622339
				11'd443: d_out <= 32'b00000000000000001001111110010110; // d_in = 1.865234, d_out = 0.623387
				11'd444: d_out <= 32'b00000000000000001001111111011011; // d_in = 1.867188, d_out = 0.624433
				11'd445: d_out <= 32'b00000000000000001010000000011111; // d_in = 1.869141, d_out = 0.625479
				11'd446: d_out <= 32'b00000000000000001010000001100100; // d_in = 1.871094, d_out = 0.626523
				11'd447: d_out <= 32'b00000000000000001010000010101000; // d_in = 1.873047, d_out = 0.627566
				11'd448: d_out <= 32'b00000000000000001010000011101100; // d_in = 1.875000, d_out = 0.628609
				11'd449: d_out <= 32'b00000000000000001010000100110001; // d_in = 1.876953, d_out = 0.629650
				11'd450: d_out <= 32'b00000000000000001010000101110101; // d_in = 1.878906, d_out = 0.630690
				11'd451: d_out <= 32'b00000000000000001010000110111001; // d_in = 1.880859, d_out = 0.631729
				11'd452: d_out <= 32'b00000000000000001010000111111101; // d_in = 1.882812, d_out = 0.632767
				11'd453: d_out <= 32'b00000000000000001010001001000001; // d_in = 1.884766, d_out = 0.633803
				11'd454: d_out <= 32'b00000000000000001010001010000101; // d_in = 1.886719, d_out = 0.634839
				11'd455: d_out <= 32'b00000000000000001010001011001001; // d_in = 1.888672, d_out = 0.635874
				11'd456: d_out <= 32'b00000000000000001010001100001100; // d_in = 1.890625, d_out = 0.636907
				11'd457: d_out <= 32'b00000000000000001010001101010000; // d_in = 1.892578, d_out = 0.637940
				11'd458: d_out <= 32'b00000000000000001010001110010100; // d_in = 1.894531, d_out = 0.638971
				11'd459: d_out <= 32'b00000000000000001010001111010111; // d_in = 1.896484, d_out = 0.640002
				11'd460: d_out <= 32'b00000000000000001010010000011011; // d_in = 1.898438, d_out = 0.641031
				11'd461: d_out <= 32'b00000000000000001010010001011110; // d_in = 1.900391, d_out = 0.642059
				11'd462: d_out <= 32'b00000000000000001010010010100001; // d_in = 1.902344, d_out = 0.643087
				11'd463: d_out <= 32'b00000000000000001010010011100101; // d_in = 1.904297, d_out = 0.644113
				11'd464: d_out <= 32'b00000000000000001010010100101000; // d_in = 1.906250, d_out = 0.645138
				11'd465: d_out <= 32'b00000000000000001010010101101011; // d_in = 1.908203, d_out = 0.646162
				11'd466: d_out <= 32'b00000000000000001010010110101110; // d_in = 1.910156, d_out = 0.647185
				11'd467: d_out <= 32'b00000000000000001010010111110001; // d_in = 1.912109, d_out = 0.648207
				11'd468: d_out <= 32'b00000000000000001010011000110100; // d_in = 1.914062, d_out = 0.649228
				11'd469: d_out <= 32'b00000000000000001010011001110111; // d_in = 1.916016, d_out = 0.650248
				11'd470: d_out <= 32'b00000000000000001010011010111001; // d_in = 1.917969, d_out = 0.651267
				11'd471: d_out <= 32'b00000000000000001010011011111100; // d_in = 1.919922, d_out = 0.652284
				11'd472: d_out <= 32'b00000000000000001010011100111111; // d_in = 1.921875, d_out = 0.653301
				11'd473: d_out <= 32'b00000000000000001010011110000001; // d_in = 1.923828, d_out = 0.654317
				11'd474: d_out <= 32'b00000000000000001010011111000100; // d_in = 1.925781, d_out = 0.655332
				11'd475: d_out <= 32'b00000000000000001010100000000110; // d_in = 1.927734, d_out = 0.656345
				11'd476: d_out <= 32'b00000000000000001010100001001001; // d_in = 1.929688, d_out = 0.657358
				11'd477: d_out <= 32'b00000000000000001010100010001011; // d_in = 1.931641, d_out = 0.658370
				11'd478: d_out <= 32'b00000000000000001010100011001101; // d_in = 1.933594, d_out = 0.659380
				11'd479: d_out <= 32'b00000000000000001010100100001111; // d_in = 1.935547, d_out = 0.660390
				11'd480: d_out <= 32'b00000000000000001010100101010001; // d_in = 1.937500, d_out = 0.661398
				11'd481: d_out <= 32'b00000000000000001010100110010011; // d_in = 1.939453, d_out = 0.662406
				11'd482: d_out <= 32'b00000000000000001010100111010101; // d_in = 1.941406, d_out = 0.663413
				11'd483: d_out <= 32'b00000000000000001010101000010111; // d_in = 1.943359, d_out = 0.664418
				11'd484: d_out <= 32'b00000000000000001010101001011001; // d_in = 1.945312, d_out = 0.665423
				11'd485: d_out <= 32'b00000000000000001010101010011011; // d_in = 1.947266, d_out = 0.666426
				11'd486: d_out <= 32'b00000000000000001010101011011101; // d_in = 1.949219, d_out = 0.667429
				11'd487: d_out <= 32'b00000000000000001010101100011110; // d_in = 1.951172, d_out = 0.668430
				11'd488: d_out <= 32'b00000000000000001010101101100000; // d_in = 1.953125, d_out = 0.669431
				11'd489: d_out <= 32'b00000000000000001010101110100001; // d_in = 1.955078, d_out = 0.670430
				11'd490: d_out <= 32'b00000000000000001010101111100011; // d_in = 1.957031, d_out = 0.671429
				11'd491: d_out <= 32'b00000000000000001010110000100100; // d_in = 1.958984, d_out = 0.672426
				11'd492: d_out <= 32'b00000000000000001010110001100101; // d_in = 1.960938, d_out = 0.673423
				11'd493: d_out <= 32'b00000000000000001010110010100111; // d_in = 1.962891, d_out = 0.674418
				11'd494: d_out <= 32'b00000000000000001010110011101000; // d_in = 1.964844, d_out = 0.675413
				11'd495: d_out <= 32'b00000000000000001010110100101001; // d_in = 1.966797, d_out = 0.676406
				11'd496: d_out <= 32'b00000000000000001010110101101010; // d_in = 1.968750, d_out = 0.677399
				11'd497: d_out <= 32'b00000000000000001010110110101011; // d_in = 1.970703, d_out = 0.678390
				11'd498: d_out <= 32'b00000000000000001010110111101100; // d_in = 1.972656, d_out = 0.679381
				11'd499: d_out <= 32'b00000000000000001010111000101101; // d_in = 1.974609, d_out = 0.680371
				11'd500: d_out <= 32'b00000000000000001010111001101110; // d_in = 1.976562, d_out = 0.681359
				11'd501: d_out <= 32'b00000000000000001010111010101110; // d_in = 1.978516, d_out = 0.682347
				11'd502: d_out <= 32'b00000000000000001010111011101111; // d_in = 1.980469, d_out = 0.683334
				11'd503: d_out <= 32'b00000000000000001010111100110000; // d_in = 1.982422, d_out = 0.684319
				11'd504: d_out <= 32'b00000000000000001010111101110000; // d_in = 1.984375, d_out = 0.685304
				11'd505: d_out <= 32'b00000000000000001010111110110001; // d_in = 1.986328, d_out = 0.686288
				11'd506: d_out <= 32'b00000000000000001010111111110001; // d_in = 1.988281, d_out = 0.687271
				11'd507: d_out <= 32'b00000000000000001011000000110001; // d_in = 1.990234, d_out = 0.688252
				11'd508: d_out <= 32'b00000000000000001011000001110010; // d_in = 1.992188, d_out = 0.689233
				11'd509: d_out <= 32'b00000000000000001011000010110010; // d_in = 1.994141, d_out = 0.690213
				11'd510: d_out <= 32'b00000000000000001011000011110010; // d_in = 1.996094, d_out = 0.691192
				11'd511: d_out <= 32'b00000000000000001011000100110010; // d_in = 1.998047, d_out = 0.692170
				11'd512: d_out <= 32'b00000000000000001011000101110010; // d_in = 2.000000, d_out = 0.693147
				11'd513: d_out <= 32'b00000000000000001011000110110010; // d_in = 2.001953, d_out = 0.694123
				11'd514: d_out <= 32'b00000000000000001011000111110010; // d_in = 2.003906, d_out = 0.695098
				11'd515: d_out <= 32'b00000000000000001011001000110010; // d_in = 2.005859, d_out = 0.696073
				11'd516: d_out <= 32'b00000000000000001011001001110010; // d_in = 2.007812, d_out = 0.697046
				11'd517: d_out <= 32'b00000000000000001011001010110001; // d_in = 2.009766, d_out = 0.698018
				11'd518: d_out <= 32'b00000000000000001011001011110001; // d_in = 2.011719, d_out = 0.698989
				11'd519: d_out <= 32'b00000000000000001011001100110001; // d_in = 2.013672, d_out = 0.699960
				11'd520: d_out <= 32'b00000000000000001011001101110000; // d_in = 2.015625, d_out = 0.700929
				11'd521: d_out <= 32'b00000000000000001011001110110000; // d_in = 2.017578, d_out = 0.701898
				11'd522: d_out <= 32'b00000000000000001011001111101111; // d_in = 2.019531, d_out = 0.702865
				11'd523: d_out <= 32'b00000000000000001011010000101110; // d_in = 2.021484, d_out = 0.703832
				11'd524: d_out <= 32'b00000000000000001011010001101110; // d_in = 2.023438, d_out = 0.704798
				11'd525: d_out <= 32'b00000000000000001011010010101101; // d_in = 2.025391, d_out = 0.705763
				11'd526: d_out <= 32'b00000000000000001011010011101100; // d_in = 2.027344, d_out = 0.706726
				11'd527: d_out <= 32'b00000000000000001011010100101011; // d_in = 2.029297, d_out = 0.707689
				11'd528: d_out <= 32'b00000000000000001011010101101010; // d_in = 2.031250, d_out = 0.708651
				11'd529: d_out <= 32'b00000000000000001011010110101001; // d_in = 2.033203, d_out = 0.709612
				11'd530: d_out <= 32'b00000000000000001011010111101000; // d_in = 2.035156, d_out = 0.710573
				11'd531: d_out <= 32'b00000000000000001011011000100111; // d_in = 2.037109, d_out = 0.711532
				11'd532: d_out <= 32'b00000000000000001011011001100110; // d_in = 2.039062, d_out = 0.712490
				11'd533: d_out <= 32'b00000000000000001011011010100100; // d_in = 2.041016, d_out = 0.713448
				11'd534: d_out <= 32'b00000000000000001011011011100011; // d_in = 2.042969, d_out = 0.714404
				11'd535: d_out <= 32'b00000000000000001011011100100010; // d_in = 2.044922, d_out = 0.715360
				11'd536: d_out <= 32'b00000000000000001011011101100000; // d_in = 2.046875, d_out = 0.716314
				11'd537: d_out <= 32'b00000000000000001011011110011111; // d_in = 2.048828, d_out = 0.717268
				11'd538: d_out <= 32'b00000000000000001011011111011101; // d_in = 2.050781, d_out = 0.718221
				11'd539: d_out <= 32'b00000000000000001011100000011100; // d_in = 2.052734, d_out = 0.719173
				11'd540: d_out <= 32'b00000000000000001011100001011010; // d_in = 2.054688, d_out = 0.720124
				11'd541: d_out <= 32'b00000000000000001011100010011000; // d_in = 2.056641, d_out = 0.721074
				11'd542: d_out <= 32'b00000000000000001011100011010111; // d_in = 2.058594, d_out = 0.722023
				11'd543: d_out <= 32'b00000000000000001011100100010101; // d_in = 2.060547, d_out = 0.722971
				11'd544: d_out <= 32'b00000000000000001011100101010011; // d_in = 2.062500, d_out = 0.723919
				11'd545: d_out <= 32'b00000000000000001011100110010001; // d_in = 2.064453, d_out = 0.724865
				11'd546: d_out <= 32'b00000000000000001011100111001111; // d_in = 2.066406, d_out = 0.725811
				11'd547: d_out <= 32'b00000000000000001011101000001101; // d_in = 2.068359, d_out = 0.726756
				11'd548: d_out <= 32'b00000000000000001011101001001011; // d_in = 2.070312, d_out = 0.727700
				11'd549: d_out <= 32'b00000000000000001011101010001000; // d_in = 2.072266, d_out = 0.728643
				11'd550: d_out <= 32'b00000000000000001011101011000110; // d_in = 2.074219, d_out = 0.729585
				11'd551: d_out <= 32'b00000000000000001011101100000100; // d_in = 2.076172, d_out = 0.730526
				11'd552: d_out <= 32'b00000000000000001011101101000001; // d_in = 2.078125, d_out = 0.731466
				11'd553: d_out <= 32'b00000000000000001011101101111111; // d_in = 2.080078, d_out = 0.732405
				11'd554: d_out <= 32'b00000000000000001011101110111100; // d_in = 2.082031, d_out = 0.733344
				11'd555: d_out <= 32'b00000000000000001011101111111010; // d_in = 2.083984, d_out = 0.734282
				11'd556: d_out <= 32'b00000000000000001011110000110111; // d_in = 2.085938, d_out = 0.735218
				11'd557: d_out <= 32'b00000000000000001011110001110101; // d_in = 2.087891, d_out = 0.736154
				11'd558: d_out <= 32'b00000000000000001011110010110010; // d_in = 2.089844, d_out = 0.737089
				11'd559: d_out <= 32'b00000000000000001011110011101111; // d_in = 2.091797, d_out = 0.738023
				11'd560: d_out <= 32'b00000000000000001011110100101100; // d_in = 2.093750, d_out = 0.738957
				11'd561: d_out <= 32'b00000000000000001011110101101001; // d_in = 2.095703, d_out = 0.739889
				11'd562: d_out <= 32'b00000000000000001011110110100110; // d_in = 2.097656, d_out = 0.740821
				11'd563: d_out <= 32'b00000000000000001011110111100011; // d_in = 2.099609, d_out = 0.741751
				11'd564: d_out <= 32'b00000000000000001011111000100000; // d_in = 2.101562, d_out = 0.742681
				11'd565: d_out <= 32'b00000000000000001011111001011101; // d_in = 2.103516, d_out = 0.743610
				11'd566: d_out <= 32'b00000000000000001011111010011010; // d_in = 2.105469, d_out = 0.744538
				11'd567: d_out <= 32'b00000000000000001011111011010111; // d_in = 2.107422, d_out = 0.745465
				11'd568: d_out <= 32'b00000000000000001011111100010100; // d_in = 2.109375, d_out = 0.746392
				11'd569: d_out <= 32'b00000000000000001011111101010000; // d_in = 2.111328, d_out = 0.747317
				11'd570: d_out <= 32'b00000000000000001011111110001101; // d_in = 2.113281, d_out = 0.748242
				11'd571: d_out <= 32'b00000000000000001011111111001001; // d_in = 2.115234, d_out = 0.749166
				11'd572: d_out <= 32'b00000000000000001100000000000110; // d_in = 2.117188, d_out = 0.750089
				11'd573: d_out <= 32'b00000000000000001100000001000010; // d_in = 2.119141, d_out = 0.751011
				11'd574: d_out <= 32'b00000000000000001100000001111111; // d_in = 2.121094, d_out = 0.751932
				11'd575: d_out <= 32'b00000000000000001100000010111011; // d_in = 2.123047, d_out = 0.752852
				11'd576: d_out <= 32'b00000000000000001100000011110111; // d_in = 2.125000, d_out = 0.753772
				11'd577: d_out <= 32'b00000000000000001100000100110011; // d_in = 2.126953, d_out = 0.754690
				11'd578: d_out <= 32'b00000000000000001100000101110000; // d_in = 2.128906, d_out = 0.755608
				11'd579: d_out <= 32'b00000000000000001100000110101100; // d_in = 2.130859, d_out = 0.756525
				11'd580: d_out <= 32'b00000000000000001100000111101000; // d_in = 2.132812, d_out = 0.757442
				11'd581: d_out <= 32'b00000000000000001100001000100100; // d_in = 2.134766, d_out = 0.758357
				11'd582: d_out <= 32'b00000000000000001100001001100000; // d_in = 2.136719, d_out = 0.759271
				11'd583: d_out <= 32'b00000000000000001100001010011011; // d_in = 2.138672, d_out = 0.760185
				11'd584: d_out <= 32'b00000000000000001100001011010111; // d_in = 2.140625, d_out = 0.761098
				11'd585: d_out <= 32'b00000000000000001100001100010011; // d_in = 2.142578, d_out = 0.762010
				11'd586: d_out <= 32'b00000000000000001100001101001111; // d_in = 2.144531, d_out = 0.762921
				11'd587: d_out <= 32'b00000000000000001100001110001010; // d_in = 2.146484, d_out = 0.763831
				11'd588: d_out <= 32'b00000000000000001100001111000110; // d_in = 2.148438, d_out = 0.764741
				11'd589: d_out <= 32'b00000000000000001100010000000010; // d_in = 2.150391, d_out = 0.765650
				11'd590: d_out <= 32'b00000000000000001100010000111101; // d_in = 2.152344, d_out = 0.766557
				11'd591: d_out <= 32'b00000000000000001100010001111001; // d_in = 2.154297, d_out = 0.767464
				11'd592: d_out <= 32'b00000000000000001100010010110100; // d_in = 2.156250, d_out = 0.768371
				11'd593: d_out <= 32'b00000000000000001100010011101111; // d_in = 2.158203, d_out = 0.769276
				11'd594: d_out <= 32'b00000000000000001100010100101011; // d_in = 2.160156, d_out = 0.770181
				11'd595: d_out <= 32'b00000000000000001100010101100110; // d_in = 2.162109, d_out = 0.771084
				11'd596: d_out <= 32'b00000000000000001100010110100001; // d_in = 2.164062, d_out = 0.771987
				11'd597: d_out <= 32'b00000000000000001100010111011100; // d_in = 2.166016, d_out = 0.772889
				11'd598: d_out <= 32'b00000000000000001100011000010111; // d_in = 2.167969, d_out = 0.773791
				11'd599: d_out <= 32'b00000000000000001100011001010010; // d_in = 2.169922, d_out = 0.774691
				11'd600: d_out <= 32'b00000000000000001100011010001101; // d_in = 2.171875, d_out = 0.775591
				11'd601: d_out <= 32'b00000000000000001100011011001000; // d_in = 2.173828, d_out = 0.776490
				11'd602: d_out <= 32'b00000000000000001100011100000011; // d_in = 2.175781, d_out = 0.777388
				11'd603: d_out <= 32'b00000000000000001100011100111110; // d_in = 2.177734, d_out = 0.778285
				11'd604: d_out <= 32'b00000000000000001100011101111000; // d_in = 2.179688, d_out = 0.779182
				11'd605: d_out <= 32'b00000000000000001100011110110011; // d_in = 2.181641, d_out = 0.780077
				11'd606: d_out <= 32'b00000000000000001100011111101110; // d_in = 2.183594, d_out = 0.780972
				11'd607: d_out <= 32'b00000000000000001100100000101000; // d_in = 2.185547, d_out = 0.781866
				11'd608: d_out <= 32'b00000000000000001100100001100011; // d_in = 2.187500, d_out = 0.782759
				11'd609: d_out <= 32'b00000000000000001100100010011101; // d_in = 2.189453, d_out = 0.783652
				11'd610: d_out <= 32'b00000000000000001100100011011000; // d_in = 2.191406, d_out = 0.784543
				11'd611: d_out <= 32'b00000000000000001100100100010010; // d_in = 2.193359, d_out = 0.785434
				11'd612: d_out <= 32'b00000000000000001100100101001101; // d_in = 2.195312, d_out = 0.786324
				11'd613: d_out <= 32'b00000000000000001100100110000111; // d_in = 2.197266, d_out = 0.787214
				11'd614: d_out <= 32'b00000000000000001100100111000001; // d_in = 2.199219, d_out = 0.788102
				11'd615: d_out <= 32'b00000000000000001100100111111011; // d_in = 2.201172, d_out = 0.788990
				11'd616: d_out <= 32'b00000000000000001100101000110101; // d_in = 2.203125, d_out = 0.789877
				11'd617: d_out <= 32'b00000000000000001100101001101111; // d_in = 2.205078, d_out = 0.790763
				11'd618: d_out <= 32'b00000000000000001100101010101001; // d_in = 2.207031, d_out = 0.791648
				11'd619: d_out <= 32'b00000000000000001100101011100011; // d_in = 2.208984, d_out = 0.792533
				11'd620: d_out <= 32'b00000000000000001100101100011101; // d_in = 2.210938, d_out = 0.793417
				11'd621: d_out <= 32'b00000000000000001100101101010111; // d_in = 2.212891, d_out = 0.794300
				11'd622: d_out <= 32'b00000000000000001100101110010001; // d_in = 2.214844, d_out = 0.795182
				11'd623: d_out <= 32'b00000000000000001100101111001011; // d_in = 2.216797, d_out = 0.796063
				11'd624: d_out <= 32'b00000000000000001100110000000101; // d_in = 2.218750, d_out = 0.796944
				11'd625: d_out <= 32'b00000000000000001100110000111110; // d_in = 2.220703, d_out = 0.797824
				11'd626: d_out <= 32'b00000000000000001100110001111000; // d_in = 2.222656, d_out = 0.798703
				11'd627: d_out <= 32'b00000000000000001100110010110001; // d_in = 2.224609, d_out = 0.799581
				11'd628: d_out <= 32'b00000000000000001100110011101011; // d_in = 2.226562, d_out = 0.800459
				11'd629: d_out <= 32'b00000000000000001100110100100100; // d_in = 2.228516, d_out = 0.801336
				11'd630: d_out <= 32'b00000000000000001100110101011110; // d_in = 2.230469, d_out = 0.802212
				11'd631: d_out <= 32'b00000000000000001100110110010111; // d_in = 2.232422, d_out = 0.803087
				11'd632: d_out <= 32'b00000000000000001100110111010000; // d_in = 2.234375, d_out = 0.803962
				11'd633: d_out <= 32'b00000000000000001100111000001010; // d_in = 2.236328, d_out = 0.804835
				11'd634: d_out <= 32'b00000000000000001100111001000011; // d_in = 2.238281, d_out = 0.805708
				11'd635: d_out <= 32'b00000000000000001100111001111100; // d_in = 2.240234, d_out = 0.806580
				11'd636: d_out <= 32'b00000000000000001100111010110101; // d_in = 2.242188, d_out = 0.807452
				11'd637: d_out <= 32'b00000000000000001100111011101110; // d_in = 2.244141, d_out = 0.808323
				11'd638: d_out <= 32'b00000000000000001100111100100111; // d_in = 2.246094, d_out = 0.809193
				11'd639: d_out <= 32'b00000000000000001100111101100000; // d_in = 2.248047, d_out = 0.810062
				11'd640: d_out <= 32'b00000000000000001100111110011001; // d_in = 2.250000, d_out = 0.810930
				11'd641: d_out <= 32'b00000000000000001100111111010010; // d_in = 2.251953, d_out = 0.811798
				11'd642: d_out <= 32'b00000000000000001101000000001011; // d_in = 2.253906, d_out = 0.812665
				11'd643: d_out <= 32'b00000000000000001101000001000100; // d_in = 2.255859, d_out = 0.813531
				11'd644: d_out <= 32'b00000000000000001101000001111100; // d_in = 2.257812, d_out = 0.814396
				11'd645: d_out <= 32'b00000000000000001101000010110101; // d_in = 2.259766, d_out = 0.815261
				11'd646: d_out <= 32'b00000000000000001101000011101110; // d_in = 2.261719, d_out = 0.816125
				11'd647: d_out <= 32'b00000000000000001101000100100110; // d_in = 2.263672, d_out = 0.816988
				11'd648: d_out <= 32'b00000000000000001101000101011111; // d_in = 2.265625, d_out = 0.817851
				11'd649: d_out <= 32'b00000000000000001101000110010111; // d_in = 2.267578, d_out = 0.818712
				11'd650: d_out <= 32'b00000000000000001101000111010000; // d_in = 2.269531, d_out = 0.819573
				11'd651: d_out <= 32'b00000000000000001101001000001000; // d_in = 2.271484, d_out = 0.820434
				11'd652: d_out <= 32'b00000000000000001101001001000000; // d_in = 2.273438, d_out = 0.821293
				11'd653: d_out <= 32'b00000000000000001101001001111001; // d_in = 2.275391, d_out = 0.822152
				11'd654: d_out <= 32'b00000000000000001101001010110001; // d_in = 2.277344, d_out = 0.823010
				11'd655: d_out <= 32'b00000000000000001101001011101001; // d_in = 2.279297, d_out = 0.823867
				11'd656: d_out <= 32'b00000000000000001101001100100001; // d_in = 2.281250, d_out = 0.824724
				11'd657: d_out <= 32'b00000000000000001101001101011001; // d_in = 2.283203, d_out = 0.825579
				11'd658: d_out <= 32'b00000000000000001101001110010001; // d_in = 2.285156, d_out = 0.826434
				11'd659: d_out <= 32'b00000000000000001101001111001001; // d_in = 2.287109, d_out = 0.827289
				11'd660: d_out <= 32'b00000000000000001101010000000001; // d_in = 2.289062, d_out = 0.828142
				11'd661: d_out <= 32'b00000000000000001101010000111001; // d_in = 2.291016, d_out = 0.828995
				11'd662: d_out <= 32'b00000000000000001101010001110001; // d_in = 2.292969, d_out = 0.829847
				11'd663: d_out <= 32'b00000000000000001101010010101001; // d_in = 2.294922, d_out = 0.830699
				11'd664: d_out <= 32'b00000000000000001101010011100000; // d_in = 2.296875, d_out = 0.831550
				11'd665: d_out <= 32'b00000000000000001101010100011000; // d_in = 2.298828, d_out = 0.832399
				11'd666: d_out <= 32'b00000000000000001101010101010000; // d_in = 2.300781, d_out = 0.833249
				11'd667: d_out <= 32'b00000000000000001101010110000111; // d_in = 2.302734, d_out = 0.834097
				11'd668: d_out <= 32'b00000000000000001101010110111111; // d_in = 2.304688, d_out = 0.834945
				11'd669: d_out <= 32'b00000000000000001101010111110110; // d_in = 2.306641, d_out = 0.835792
				11'd670: d_out <= 32'b00000000000000001101011000101110; // d_in = 2.308594, d_out = 0.836639
				11'd671: d_out <= 32'b00000000000000001101011001100101; // d_in = 2.310547, d_out = 0.837484
				11'd672: d_out <= 32'b00000000000000001101011010011101; // d_in = 2.312500, d_out = 0.838329
				11'd673: d_out <= 32'b00000000000000001101011011010100; // d_in = 2.314453, d_out = 0.839173
				11'd674: d_out <= 32'b00000000000000001101011100001011; // d_in = 2.316406, d_out = 0.840017
				11'd675: d_out <= 32'b00000000000000001101011101000011; // d_in = 2.318359, d_out = 0.840860
				11'd676: d_out <= 32'b00000000000000001101011101111010; // d_in = 2.320312, d_out = 0.841702
				11'd677: d_out <= 32'b00000000000000001101011110110001; // d_in = 2.322266, d_out = 0.842543
				11'd678: d_out <= 32'b00000000000000001101011111101000; // d_in = 2.324219, d_out = 0.843384
				11'd679: d_out <= 32'b00000000000000001101100000011111; // d_in = 2.326172, d_out = 0.844224
				11'd680: d_out <= 32'b00000000000000001101100001010110; // d_in = 2.328125, d_out = 0.845063
				11'd681: d_out <= 32'b00000000000000001101100010001101; // d_in = 2.330078, d_out = 0.845902
				11'd682: d_out <= 32'b00000000000000001101100011000100; // d_in = 2.332031, d_out = 0.846740
				11'd683: d_out <= 32'b00000000000000001101100011111011; // d_in = 2.333984, d_out = 0.847577
				11'd684: d_out <= 32'b00000000000000001101100100110010; // d_in = 2.335938, d_out = 0.848413
				11'd685: d_out <= 32'b00000000000000001101100101101000; // d_in = 2.337891, d_out = 0.849249
				11'd686: d_out <= 32'b00000000000000001101100110011111; // d_in = 2.339844, d_out = 0.850084
				11'd687: d_out <= 32'b00000000000000001101100111010110; // d_in = 2.341797, d_out = 0.850919
				11'd688: d_out <= 32'b00000000000000001101101000001100; // d_in = 2.343750, d_out = 0.851752
				11'd689: d_out <= 32'b00000000000000001101101001000011; // d_in = 2.345703, d_out = 0.852585
				11'd690: d_out <= 32'b00000000000000001101101001111010; // d_in = 2.347656, d_out = 0.853417
				11'd691: d_out <= 32'b00000000000000001101101010110000; // d_in = 2.349609, d_out = 0.854249
				11'd692: d_out <= 32'b00000000000000001101101011100111; // d_in = 2.351562, d_out = 0.855080
				11'd693: d_out <= 32'b00000000000000001101101100011101; // d_in = 2.353516, d_out = 0.855910
				11'd694: d_out <= 32'b00000000000000001101101101010011; // d_in = 2.355469, d_out = 0.856740
				11'd695: d_out <= 32'b00000000000000001101101110001010; // d_in = 2.357422, d_out = 0.857569
				11'd696: d_out <= 32'b00000000000000001101101111000000; // d_in = 2.359375, d_out = 0.858397
				11'd697: d_out <= 32'b00000000000000001101101111110110; // d_in = 2.361328, d_out = 0.859224
				11'd698: d_out <= 32'b00000000000000001101110000101100; // d_in = 2.363281, d_out = 0.860051
				11'd699: d_out <= 32'b00000000000000001101110001100010; // d_in = 2.365234, d_out = 0.860877
				11'd700: d_out <= 32'b00000000000000001101110010011001; // d_in = 2.367188, d_out = 0.861703
				11'd701: d_out <= 32'b00000000000000001101110011001111; // d_in = 2.369141, d_out = 0.862527
				11'd702: d_out <= 32'b00000000000000001101110100000101; // d_in = 2.371094, d_out = 0.863351
				11'd703: d_out <= 32'b00000000000000001101110100111011; // d_in = 2.373047, d_out = 0.864175
				11'd704: d_out <= 32'b00000000000000001101110101110000; // d_in = 2.375000, d_out = 0.864997
				11'd705: d_out <= 32'b00000000000000001101110110100110; // d_in = 2.376953, d_out = 0.865819
				11'd706: d_out <= 32'b00000000000000001101110111011100; // d_in = 2.378906, d_out = 0.866641
				11'd707: d_out <= 32'b00000000000000001101111000010010; // d_in = 2.380859, d_out = 0.867462
				11'd708: d_out <= 32'b00000000000000001101111001001000; // d_in = 2.382812, d_out = 0.868282
				11'd709: d_out <= 32'b00000000000000001101111001111101; // d_in = 2.384766, d_out = 0.869101
				11'd710: d_out <= 32'b00000000000000001101111010110011; // d_in = 2.386719, d_out = 0.869920
				11'd711: d_out <= 32'b00000000000000001101111011101001; // d_in = 2.388672, d_out = 0.870738
				11'd712: d_out <= 32'b00000000000000001101111100011110; // d_in = 2.390625, d_out = 0.871555
				11'd713: d_out <= 32'b00000000000000001101111101010100; // d_in = 2.392578, d_out = 0.872371
				11'd714: d_out <= 32'b00000000000000001101111110001001; // d_in = 2.394531, d_out = 0.873187
				11'd715: d_out <= 32'b00000000000000001101111110111111; // d_in = 2.396484, d_out = 0.874003
				11'd716: d_out <= 32'b00000000000000001101111111110100; // d_in = 2.398438, d_out = 0.874817
				11'd717: d_out <= 32'b00000000000000001110000000101001; // d_in = 2.400391, d_out = 0.875631
				11'd718: d_out <= 32'b00000000000000001110000001011111; // d_in = 2.402344, d_out = 0.876445
				11'd719: d_out <= 32'b00000000000000001110000010010100; // d_in = 2.404297, d_out = 0.877258
				11'd720: d_out <= 32'b00000000000000001110000011001001; // d_in = 2.406250, d_out = 0.878070
				11'd721: d_out <= 32'b00000000000000001110000011111110; // d_in = 2.408203, d_out = 0.878881
				11'd722: d_out <= 32'b00000000000000001110000100110011; // d_in = 2.410156, d_out = 0.879692
				11'd723: d_out <= 32'b00000000000000001110000101101001; // d_in = 2.412109, d_out = 0.880502
				11'd724: d_out <= 32'b00000000000000001110000110011110; // d_in = 2.414062, d_out = 0.881311
				11'd725: d_out <= 32'b00000000000000001110000111010011; // d_in = 2.416016, d_out = 0.882120
				11'd726: d_out <= 32'b00000000000000001110001000001000; // d_in = 2.417969, d_out = 0.882928
				11'd727: d_out <= 32'b00000000000000001110001000111100; // d_in = 2.419922, d_out = 0.883735
				11'd728: d_out <= 32'b00000000000000001110001001110001; // d_in = 2.421875, d_out = 0.884542
				11'd729: d_out <= 32'b00000000000000001110001010100110; // d_in = 2.423828, d_out = 0.885348
				11'd730: d_out <= 32'b00000000000000001110001011011011; // d_in = 2.425781, d_out = 0.886154
				11'd731: d_out <= 32'b00000000000000001110001100010000; // d_in = 2.427734, d_out = 0.886958
				11'd732: d_out <= 32'b00000000000000001110001101000100; // d_in = 2.429688, d_out = 0.887763
				11'd733: d_out <= 32'b00000000000000001110001101111001; // d_in = 2.431641, d_out = 0.888566
				11'd734: d_out <= 32'b00000000000000001110001110101110; // d_in = 2.433594, d_out = 0.889369
				11'd735: d_out <= 32'b00000000000000001110001111100010; // d_in = 2.435547, d_out = 0.890171
				11'd736: d_out <= 32'b00000000000000001110010000010111; // d_in = 2.437500, d_out = 0.890973
				11'd737: d_out <= 32'b00000000000000001110010001001011; // d_in = 2.439453, d_out = 0.891774
				11'd738: d_out <= 32'b00000000000000001110010010000000; // d_in = 2.441406, d_out = 0.892574
				11'd739: d_out <= 32'b00000000000000001110010010110100; // d_in = 2.443359, d_out = 0.893374
				11'd740: d_out <= 32'b00000000000000001110010011101001; // d_in = 2.445312, d_out = 0.894173
				11'd741: d_out <= 32'b00000000000000001110010100011101; // d_in = 2.447266, d_out = 0.894971
				11'd742: d_out <= 32'b00000000000000001110010101010001; // d_in = 2.449219, d_out = 0.895769
				11'd743: d_out <= 32'b00000000000000001110010110000101; // d_in = 2.451172, d_out = 0.896566
				11'd744: d_out <= 32'b00000000000000001110010110111010; // d_in = 2.453125, d_out = 0.897363
				11'd745: d_out <= 32'b00000000000000001110010111101110; // d_in = 2.455078, d_out = 0.898159
				11'd746: d_out <= 32'b00000000000000001110011000100010; // d_in = 2.457031, d_out = 0.898954
				11'd747: d_out <= 32'b00000000000000001110011001010110; // d_in = 2.458984, d_out = 0.899748
				11'd748: d_out <= 32'b00000000000000001110011010001010; // d_in = 2.460938, d_out = 0.900542
				11'd749: d_out <= 32'b00000000000000001110011010111110; // d_in = 2.462891, d_out = 0.901336
				11'd750: d_out <= 32'b00000000000000001110011011110010; // d_in = 2.464844, d_out = 0.902128
				11'd751: d_out <= 32'b00000000000000001110011100100110; // d_in = 2.466797, d_out = 0.902920
				11'd752: d_out <= 32'b00000000000000001110011101011010; // d_in = 2.468750, d_out = 0.903712
				11'd753: d_out <= 32'b00000000000000001110011110001101; // d_in = 2.470703, d_out = 0.904503
				11'd754: d_out <= 32'b00000000000000001110011111000001; // d_in = 2.472656, d_out = 0.905293
				11'd755: d_out <= 32'b00000000000000001110011111110101; // d_in = 2.474609, d_out = 0.906083
				11'd756: d_out <= 32'b00000000000000001110100000101001; // d_in = 2.476562, d_out = 0.906872
				11'd757: d_out <= 32'b00000000000000001110100001011100; // d_in = 2.478516, d_out = 0.907660
				11'd758: d_out <= 32'b00000000000000001110100010010000; // d_in = 2.480469, d_out = 0.908448
				11'd759: d_out <= 32'b00000000000000001110100011000100; // d_in = 2.482422, d_out = 0.909235
				11'd760: d_out <= 32'b00000000000000001110100011110111; // d_in = 2.484375, d_out = 0.910021
				11'd761: d_out <= 32'b00000000000000001110100100101011; // d_in = 2.486328, d_out = 0.910807
				11'd762: d_out <= 32'b00000000000000001110100101011110; // d_in = 2.488281, d_out = 0.911592
				11'd763: d_out <= 32'b00000000000000001110100110010010; // d_in = 2.490234, d_out = 0.912377
				11'd764: d_out <= 32'b00000000000000001110100111000101; // d_in = 2.492188, d_out = 0.913161
				11'd765: d_out <= 32'b00000000000000001110100111111000; // d_in = 2.494141, d_out = 0.913944
				11'd766: d_out <= 32'b00000000000000001110101000101100; // d_in = 2.496094, d_out = 0.914727
				11'd767: d_out <= 32'b00000000000000001110101001011111; // d_in = 2.498047, d_out = 0.915509
				11'd768: d_out <= 32'b00000000000000001110101010010010; // d_in = 2.500000, d_out = 0.916291
				11'd769: d_out <= 32'b00000000000000001110101011000101; // d_in = 2.501953, d_out = 0.917072
				11'd770: d_out <= 32'b00000000000000001110101011111000; // d_in = 2.503906, d_out = 0.917852
				11'd771: d_out <= 32'b00000000000000001110101100101011; // d_in = 2.505859, d_out = 0.918632
				11'd772: d_out <= 32'b00000000000000001110101101011111; // d_in = 2.507812, d_out = 0.919411
				11'd773: d_out <= 32'b00000000000000001110101110010010; // d_in = 2.509766, d_out = 0.920189
				11'd774: d_out <= 32'b00000000000000001110101111000101; // d_in = 2.511719, d_out = 0.920967
				11'd775: d_out <= 32'b00000000000000001110101111110111; // d_in = 2.513672, d_out = 0.921745
				11'd776: d_out <= 32'b00000000000000001110110000101010; // d_in = 2.515625, d_out = 0.922521
				11'd777: d_out <= 32'b00000000000000001110110001011101; // d_in = 2.517578, d_out = 0.923297
				11'd778: d_out <= 32'b00000000000000001110110010010000; // d_in = 2.519531, d_out = 0.924073
				11'd779: d_out <= 32'b00000000000000001110110011000011; // d_in = 2.521484, d_out = 0.924848
				11'd780: d_out <= 32'b00000000000000001110110011110110; // d_in = 2.523438, d_out = 0.925622
				11'd781: d_out <= 32'b00000000000000001110110100101000; // d_in = 2.525391, d_out = 0.926396
				11'd782: d_out <= 32'b00000000000000001110110101011011; // d_in = 2.527344, d_out = 0.927169
				11'd783: d_out <= 32'b00000000000000001110110110001110; // d_in = 2.529297, d_out = 0.927941
				11'd784: d_out <= 32'b00000000000000001110110111000000; // d_in = 2.531250, d_out = 0.928713
				11'd785: d_out <= 32'b00000000000000001110110111110011; // d_in = 2.533203, d_out = 0.929485
				11'd786: d_out <= 32'b00000000000000001110111000100101; // d_in = 2.535156, d_out = 0.930255
				11'd787: d_out <= 32'b00000000000000001110111001011000; // d_in = 2.537109, d_out = 0.931025
				11'd788: d_out <= 32'b00000000000000001110111010001010; // d_in = 2.539062, d_out = 0.931795
				11'd789: d_out <= 32'b00000000000000001110111010111101; // d_in = 2.541016, d_out = 0.932564
				11'd790: d_out <= 32'b00000000000000001110111011101111; // d_in = 2.542969, d_out = 0.933332
				11'd791: d_out <= 32'b00000000000000001110111100100001; // d_in = 2.544922, d_out = 0.934100
				11'd792: d_out <= 32'b00000000000000001110111101010011; // d_in = 2.546875, d_out = 0.934867
				11'd793: d_out <= 32'b00000000000000001110111110000110; // d_in = 2.548828, d_out = 0.935634
				11'd794: d_out <= 32'b00000000000000001110111110111000; // d_in = 2.550781, d_out = 0.936400
				11'd795: d_out <= 32'b00000000000000001110111111101010; // d_in = 2.552734, d_out = 0.937165
				11'd796: d_out <= 32'b00000000000000001111000000011100; // d_in = 2.554688, d_out = 0.937930
				11'd797: d_out <= 32'b00000000000000001111000001001110; // d_in = 2.556641, d_out = 0.938694
				11'd798: d_out <= 32'b00000000000000001111000010000000; // d_in = 2.558594, d_out = 0.939458
				11'd799: d_out <= 32'b00000000000000001111000010110010; // d_in = 2.560547, d_out = 0.940221
				11'd800: d_out <= 32'b00000000000000001111000011100100; // d_in = 2.562500, d_out = 0.940983
				11'd801: d_out <= 32'b00000000000000001111000100010110; // d_in = 2.564453, d_out = 0.941745
				11'd802: d_out <= 32'b00000000000000001111000101001000; // d_in = 2.566406, d_out = 0.942507
				11'd803: d_out <= 32'b00000000000000001111000101111010; // d_in = 2.568359, d_out = 0.943267
				11'd804: d_out <= 32'b00000000000000001111000110101100; // d_in = 2.570312, d_out = 0.944027
				11'd805: d_out <= 32'b00000000000000001111000111011110; // d_in = 2.572266, d_out = 0.944787
				11'd806: d_out <= 32'b00000000000000001111001000001111; // d_in = 2.574219, d_out = 0.945546
				11'd807: d_out <= 32'b00000000000000001111001001000001; // d_in = 2.576172, d_out = 0.946305
				11'd808: d_out <= 32'b00000000000000001111001001110011; // d_in = 2.578125, d_out = 0.947062
				11'd809: d_out <= 32'b00000000000000001111001010100100; // d_in = 2.580078, d_out = 0.947820
				11'd810: d_out <= 32'b00000000000000001111001011010110; // d_in = 2.582031, d_out = 0.948576
				11'd811: d_out <= 32'b00000000000000001111001100000111; // d_in = 2.583984, d_out = 0.949333
				11'd812: d_out <= 32'b00000000000000001111001100111001; // d_in = 2.585938, d_out = 0.950088
				11'd813: d_out <= 32'b00000000000000001111001101101010; // d_in = 2.587891, d_out = 0.950843
				11'd814: d_out <= 32'b00000000000000001111001110011100; // d_in = 2.589844, d_out = 0.951598
				11'd815: d_out <= 32'b00000000000000001111001111001101; // d_in = 2.591797, d_out = 0.952351
				11'd816: d_out <= 32'b00000000000000001111001111111111; // d_in = 2.593750, d_out = 0.953105
				11'd817: d_out <= 32'b00000000000000001111010000110000; // d_in = 2.595703, d_out = 0.953857
				11'd818: d_out <= 32'b00000000000000001111010001100001; // d_in = 2.597656, d_out = 0.954610
				11'd819: d_out <= 32'b00000000000000001111010010010011; // d_in = 2.599609, d_out = 0.955361
				11'd820: d_out <= 32'b00000000000000001111010011000100; // d_in = 2.601562, d_out = 0.956112
				11'd821: d_out <= 32'b00000000000000001111010011110101; // d_in = 2.603516, d_out = 0.956863
				11'd822: d_out <= 32'b00000000000000001111010100100110; // d_in = 2.605469, d_out = 0.957613
				11'd823: d_out <= 32'b00000000000000001111010101010111; // d_in = 2.607422, d_out = 0.958362
				11'd824: d_out <= 32'b00000000000000001111010110001000; // d_in = 2.609375, d_out = 0.959111
				11'd825: d_out <= 32'b00000000000000001111010110111001; // d_in = 2.611328, d_out = 0.959859
				11'd826: d_out <= 32'b00000000000000001111010111101010; // d_in = 2.613281, d_out = 0.960607
				11'd827: d_out <= 32'b00000000000000001111011000011011; // d_in = 2.615234, d_out = 0.961354
				11'd828: d_out <= 32'b00000000000000001111011001001100; // d_in = 2.617188, d_out = 0.962100
				11'd829: d_out <= 32'b00000000000000001111011001111101; // d_in = 2.619141, d_out = 0.962846
				11'd830: d_out <= 32'b00000000000000001111011010101110; // d_in = 2.621094, d_out = 0.963592
				11'd831: d_out <= 32'b00000000000000001111011011011111; // d_in = 2.623047, d_out = 0.964337
				11'd832: d_out <= 32'b00000000000000001111011100010000; // d_in = 2.625000, d_out = 0.965081
				11'd833: d_out <= 32'b00000000000000001111011101000000; // d_in = 2.626953, d_out = 0.965825
				11'd834: d_out <= 32'b00000000000000001111011101110001; // d_in = 2.628906, d_out = 0.966568
				11'd835: d_out <= 32'b00000000000000001111011110100010; // d_in = 2.630859, d_out = 0.967311
				11'd836: d_out <= 32'b00000000000000001111011111010010; // d_in = 2.632812, d_out = 0.968053
				11'd837: d_out <= 32'b00000000000000001111100000000011; // d_in = 2.634766, d_out = 0.968794
				11'd838: d_out <= 32'b00000000000000001111100000110011; // d_in = 2.636719, d_out = 0.969535
				11'd839: d_out <= 32'b00000000000000001111100001100100; // d_in = 2.638672, d_out = 0.970276
				11'd840: d_out <= 32'b00000000000000001111100010010100; // d_in = 2.640625, d_out = 0.971016
				11'd841: d_out <= 32'b00000000000000001111100011000101; // d_in = 2.642578, d_out = 0.971755
				11'd842: d_out <= 32'b00000000000000001111100011110101; // d_in = 2.644531, d_out = 0.972494
				11'd843: d_out <= 32'b00000000000000001111100100100110; // d_in = 2.646484, d_out = 0.973232
				11'd844: d_out <= 32'b00000000000000001111100101010110; // d_in = 2.648438, d_out = 0.973970
				11'd845: d_out <= 32'b00000000000000001111100110000110; // d_in = 2.650391, d_out = 0.974707
				11'd846: d_out <= 32'b00000000000000001111100110110111; // d_in = 2.652344, d_out = 0.975444
				11'd847: d_out <= 32'b00000000000000001111100111100111; // d_in = 2.654297, d_out = 0.976180
				11'd848: d_out <= 32'b00000000000000001111101000010111; // d_in = 2.656250, d_out = 0.976915
				11'd849: d_out <= 32'b00000000000000001111101001000111; // d_in = 2.658203, d_out = 0.977650
				11'd850: d_out <= 32'b00000000000000001111101001110111; // d_in = 2.660156, d_out = 0.978385
				11'd851: d_out <= 32'b00000000000000001111101010101000; // d_in = 2.662109, d_out = 0.979119
				11'd852: d_out <= 32'b00000000000000001111101011011000; // d_in = 2.664062, d_out = 0.979852
				11'd853: d_out <= 32'b00000000000000001111101100001000; // d_in = 2.666016, d_out = 0.980585
				11'd854: d_out <= 32'b00000000000000001111101100111000; // d_in = 2.667969, d_out = 0.981317
				11'd855: d_out <= 32'b00000000000000001111101101101000; // d_in = 2.669922, d_out = 0.982049
				11'd856: d_out <= 32'b00000000000000001111101110011000; // d_in = 2.671875, d_out = 0.982780
				11'd857: d_out <= 32'b00000000000000001111101111000111; // d_in = 2.673828, d_out = 0.983511
				11'd858: d_out <= 32'b00000000000000001111101111110111; // d_in = 2.675781, d_out = 0.984241
				11'd859: d_out <= 32'b00000000000000001111110000100111; // d_in = 2.677734, d_out = 0.984971
				11'd860: d_out <= 32'b00000000000000001111110001010111; // d_in = 2.679688, d_out = 0.985700
				11'd861: d_out <= 32'b00000000000000001111110010000111; // d_in = 2.681641, d_out = 0.986429
				11'd862: d_out <= 32'b00000000000000001111110010110110; // d_in = 2.683594, d_out = 0.987157
				11'd863: d_out <= 32'b00000000000000001111110011100110; // d_in = 2.685547, d_out = 0.987884
				11'd864: d_out <= 32'b00000000000000001111110100010110; // d_in = 2.687500, d_out = 0.988611
				11'd865: d_out <= 32'b00000000000000001111110101000101; // d_in = 2.689453, d_out = 0.989338
				11'd866: d_out <= 32'b00000000000000001111110101110101; // d_in = 2.691406, d_out = 0.990064
				11'd867: d_out <= 32'b00000000000000001111110110100100; // d_in = 2.693359, d_out = 0.990789
				11'd868: d_out <= 32'b00000000000000001111110111010100; // d_in = 2.695312, d_out = 0.991514
				11'd869: d_out <= 32'b00000000000000001111111000000011; // d_in = 2.697266, d_out = 0.992239
				11'd870: d_out <= 32'b00000000000000001111111000110011; // d_in = 2.699219, d_out = 0.992962
				11'd871: d_out <= 32'b00000000000000001111111001100010; // d_in = 2.701172, d_out = 0.993686
				11'd872: d_out <= 32'b00000000000000001111111010010010; // d_in = 2.703125, d_out = 0.994409
				11'd873: d_out <= 32'b00000000000000001111111011000001; // d_in = 2.705078, d_out = 0.995131
				11'd874: d_out <= 32'b00000000000000001111111011110000; // d_in = 2.707031, d_out = 0.995853
				11'd875: d_out <= 32'b00000000000000001111111100011111; // d_in = 2.708984, d_out = 0.996574
				11'd876: d_out <= 32'b00000000000000001111111101001111; // d_in = 2.710938, d_out = 0.997295
				11'd877: d_out <= 32'b00000000000000001111111101111110; // d_in = 2.712891, d_out = 0.998015
				11'd878: d_out <= 32'b00000000000000001111111110101101; // d_in = 2.714844, d_out = 0.998734
				11'd879: d_out <= 32'b00000000000000001111111111011100; // d_in = 2.716797, d_out = 0.999454
				11'd880: d_out <= 32'b00000000000000010000000000001011; // d_in = 2.718750, d_out = 1.000172
				11'd881: d_out <= 32'b00000000000000010000000000111010; // d_in = 2.720703, d_out = 1.000890
				11'd882: d_out <= 32'b00000000000000010000000001101001; // d_in = 2.722656, d_out = 1.001608
				11'd883: d_out <= 32'b00000000000000010000000010011000; // d_in = 2.724609, d_out = 1.002325
				11'd884: d_out <= 32'b00000000000000010000000011000111; // d_in = 2.726562, d_out = 1.003042
				11'd885: d_out <= 32'b00000000000000010000000011110110; // d_in = 2.728516, d_out = 1.003758
				11'd886: d_out <= 32'b00000000000000010000000100100101; // d_in = 2.730469, d_out = 1.004473
				11'd887: d_out <= 32'b00000000000000010000000101010100; // d_in = 2.732422, d_out = 1.005188
				11'd888: d_out <= 32'b00000000000000010000000110000011; // d_in = 2.734375, d_out = 1.005903
				11'd889: d_out <= 32'b00000000000000010000000110110010; // d_in = 2.736328, d_out = 1.006617
				11'd890: d_out <= 32'b00000000000000010000000111100000; // d_in = 2.738281, d_out = 1.007330
				11'd891: d_out <= 32'b00000000000000010000001000001111; // d_in = 2.740234, d_out = 1.008043
				11'd892: d_out <= 32'b00000000000000010000001000111110; // d_in = 2.742188, d_out = 1.008756
				11'd893: d_out <= 32'b00000000000000010000001001101100; // d_in = 2.744141, d_out = 1.009468
				11'd894: d_out <= 32'b00000000000000010000001010011011; // d_in = 2.746094, d_out = 1.010179
				11'd895: d_out <= 32'b00000000000000010000001011001010; // d_in = 2.748047, d_out = 1.010890
				11'd896: d_out <= 32'b00000000000000010000001011111000; // d_in = 2.750000, d_out = 1.011601
				11'd897: d_out <= 32'b00000000000000010000001100100111; // d_in = 2.751953, d_out = 1.012311
				11'd898: d_out <= 32'b00000000000000010000001101010101; // d_in = 2.753906, d_out = 1.013020
				11'd899: d_out <= 32'b00000000000000010000001110000100; // d_in = 2.755859, d_out = 1.013729
				11'd900: d_out <= 32'b00000000000000010000001110110010; // d_in = 2.757812, d_out = 1.014438
				11'd901: d_out <= 32'b00000000000000010000001111100001; // d_in = 2.759766, d_out = 1.015146
				11'd902: d_out <= 32'b00000000000000010000010000001111; // d_in = 2.761719, d_out = 1.015853
				11'd903: d_out <= 32'b00000000000000010000010000111101; // d_in = 2.763672, d_out = 1.016560
				11'd904: d_out <= 32'b00000000000000010000010001101100; // d_in = 2.765625, d_out = 1.017267
				11'd905: d_out <= 32'b00000000000000010000010010011010; // d_in = 2.767578, d_out = 1.017973
				11'd906: d_out <= 32'b00000000000000010000010011001000; // d_in = 2.769531, d_out = 1.018678
				11'd907: d_out <= 32'b00000000000000010000010011110110; // d_in = 2.771484, d_out = 1.019383
				11'd908: d_out <= 32'b00000000000000010000010100100100; // d_in = 2.773438, d_out = 1.020088
				11'd909: d_out <= 32'b00000000000000010000010101010011; // d_in = 2.775391, d_out = 1.020792
				11'd910: d_out <= 32'b00000000000000010000010110000001; // d_in = 2.777344, d_out = 1.021495
				11'd911: d_out <= 32'b00000000000000010000010110101111; // d_in = 2.779297, d_out = 1.022198
				11'd912: d_out <= 32'b00000000000000010000010111011101; // d_in = 2.781250, d_out = 1.022900
				11'd913: d_out <= 32'b00000000000000010000011000001011; // d_in = 2.783203, d_out = 1.023602
				11'd914: d_out <= 32'b00000000000000010000011000111001; // d_in = 2.785156, d_out = 1.024304
				11'd915: d_out <= 32'b00000000000000010000011001100111; // d_in = 2.787109, d_out = 1.025005
				11'd916: d_out <= 32'b00000000000000010000011010010101; // d_in = 2.789062, d_out = 1.025706
				11'd917: d_out <= 32'b00000000000000010000011011000011; // d_in = 2.791016, d_out = 1.026406
				11'd918: d_out <= 32'b00000000000000010000011011110000; // d_in = 2.792969, d_out = 1.027105
				11'd919: d_out <= 32'b00000000000000010000011100011110; // d_in = 2.794922, d_out = 1.027804
				11'd920: d_out <= 32'b00000000000000010000011101001100; // d_in = 2.796875, d_out = 1.028503
				11'd921: d_out <= 32'b00000000000000010000011101111010; // d_in = 2.798828, d_out = 1.029201
				11'd922: d_out <= 32'b00000000000000010000011110100111; // d_in = 2.800781, d_out = 1.029898
				11'd923: d_out <= 32'b00000000000000010000011111010101; // d_in = 2.802734, d_out = 1.030596
				11'd924: d_out <= 32'b00000000000000010000100000000011; // d_in = 2.804688, d_out = 1.031292
				11'd925: d_out <= 32'b00000000000000010000100000110000; // d_in = 2.806641, d_out = 1.031988
				11'd926: d_out <= 32'b00000000000000010000100001011110; // d_in = 2.808594, d_out = 1.032684
				11'd927: d_out <= 32'b00000000000000010000100010001100; // d_in = 2.810547, d_out = 1.033379
				11'd928: d_out <= 32'b00000000000000010000100010111001; // d_in = 2.812500, d_out = 1.034074
				11'd929: d_out <= 32'b00000000000000010000100011100111; // d_in = 2.814453, d_out = 1.034768
				11'd930: d_out <= 32'b00000000000000010000100100010100; // d_in = 2.816406, d_out = 1.035462
				11'd931: d_out <= 32'b00000000000000010000100101000001; // d_in = 2.818359, d_out = 1.036155
				11'd932: d_out <= 32'b00000000000000010000100101101111; // d_in = 2.820312, d_out = 1.036848
				11'd933: d_out <= 32'b00000000000000010000100110011100; // d_in = 2.822266, d_out = 1.037540
				11'd934: d_out <= 32'b00000000000000010000100111001010; // d_in = 2.824219, d_out = 1.038232
				11'd935: d_out <= 32'b00000000000000010000100111110111; // d_in = 2.826172, d_out = 1.038923
				11'd936: d_out <= 32'b00000000000000010000101000100100; // d_in = 2.828125, d_out = 1.039614
				11'd937: d_out <= 32'b00000000000000010000101001010001; // d_in = 2.830078, d_out = 1.040304
				11'd938: d_out <= 32'b00000000000000010000101001111111; // d_in = 2.832031, d_out = 1.040994
				11'd939: d_out <= 32'b00000000000000010000101010101100; // d_in = 2.833984, d_out = 1.041684
				11'd940: d_out <= 32'b00000000000000010000101011011001; // d_in = 2.835938, d_out = 1.042373
				11'd941: d_out <= 32'b00000000000000010000101100000110; // d_in = 2.837891, d_out = 1.043061
				11'd942: d_out <= 32'b00000000000000010000101100110011; // d_in = 2.839844, d_out = 1.043749
				11'd943: d_out <= 32'b00000000000000010000101101100000; // d_in = 2.841797, d_out = 1.044437
				11'd944: d_out <= 32'b00000000000000010000101110001101; // d_in = 2.843750, d_out = 1.045124
				11'd945: d_out <= 32'b00000000000000010000101110111010; // d_in = 2.845703, d_out = 1.045810
				11'd946: d_out <= 32'b00000000000000010000101111100111; // d_in = 2.847656, d_out = 1.046496
				11'd947: d_out <= 32'b00000000000000010000110000010100; // d_in = 2.849609, d_out = 1.047182
				11'd948: d_out <= 32'b00000000000000010000110001000001; // d_in = 2.851562, d_out = 1.047867
				11'd949: d_out <= 32'b00000000000000010000110001101110; // d_in = 2.853516, d_out = 1.048552
				11'd950: d_out <= 32'b00000000000000010000110010011011; // d_in = 2.855469, d_out = 1.049236
				11'd951: d_out <= 32'b00000000000000010000110011001000; // d_in = 2.857422, d_out = 1.049920
				11'd952: d_out <= 32'b00000000000000010000110011110100; // d_in = 2.859375, d_out = 1.050603
				11'd953: d_out <= 32'b00000000000000010000110100100001; // d_in = 2.861328, d_out = 1.051286
				11'd954: d_out <= 32'b00000000000000010000110101001110; // d_in = 2.863281, d_out = 1.051968
				11'd955: d_out <= 32'b00000000000000010000110101111010; // d_in = 2.865234, d_out = 1.052650
				11'd956: d_out <= 32'b00000000000000010000110110100111; // d_in = 2.867188, d_out = 1.053332
				11'd957: d_out <= 32'b00000000000000010000110111010100; // d_in = 2.869141, d_out = 1.054013
				11'd958: d_out <= 32'b00000000000000010000111000000000; // d_in = 2.871094, d_out = 1.054693
				11'd959: d_out <= 32'b00000000000000010000111000101101; // d_in = 2.873047, d_out = 1.055373
				11'd960: d_out <= 32'b00000000000000010000111001011001; // d_in = 2.875000, d_out = 1.056053
				11'd961: d_out <= 32'b00000000000000010000111010000110; // d_in = 2.876953, d_out = 1.056732
				11'd962: d_out <= 32'b00000000000000010000111010110010; // d_in = 2.878906, d_out = 1.057410
				11'd963: d_out <= 32'b00000000000000010000111011011111; // d_in = 2.880859, d_out = 1.058089
				11'd964: d_out <= 32'b00000000000000010000111100001011; // d_in = 2.882812, d_out = 1.058766
				11'd965: d_out <= 32'b00000000000000010000111100111000; // d_in = 2.884766, d_out = 1.059444
				11'd966: d_out <= 32'b00000000000000010000111101100100; // d_in = 2.886719, d_out = 1.060120
				11'd967: d_out <= 32'b00000000000000010000111110010000; // d_in = 2.888672, d_out = 1.060797
				11'd968: d_out <= 32'b00000000000000010000111110111101; // d_in = 2.890625, d_out = 1.061473
				11'd969: d_out <= 32'b00000000000000010000111111101001; // d_in = 2.892578, d_out = 1.062148
				11'd970: d_out <= 32'b00000000000000010001000000010101; // d_in = 2.894531, d_out = 1.062823
				11'd971: d_out <= 32'b00000000000000010001000001000001; // d_in = 2.896484, d_out = 1.063498
				11'd972: d_out <= 32'b00000000000000010001000001101110; // d_in = 2.898438, d_out = 1.064172
				11'd973: d_out <= 32'b00000000000000010001000010011010; // d_in = 2.900391, d_out = 1.064845
				11'd974: d_out <= 32'b00000000000000010001000011000110; // d_in = 2.902344, d_out = 1.065519
				11'd975: d_out <= 32'b00000000000000010001000011110010; // d_in = 2.904297, d_out = 1.066191
				11'd976: d_out <= 32'b00000000000000010001000100011110; // d_in = 2.906250, d_out = 1.066864
				11'd977: d_out <= 32'b00000000000000010001000101001010; // d_in = 2.908203, d_out = 1.067535
				11'd978: d_out <= 32'b00000000000000010001000101110110; // d_in = 2.910156, d_out = 1.068207
				11'd979: d_out <= 32'b00000000000000010001000110100010; // d_in = 2.912109, d_out = 1.068878
				11'd980: d_out <= 32'b00000000000000010001000111001110; // d_in = 2.914062, d_out = 1.069548
				11'd981: d_out <= 32'b00000000000000010001000111111010; // d_in = 2.916016, d_out = 1.070218
				11'd982: d_out <= 32'b00000000000000010001001000100110; // d_in = 2.917969, d_out = 1.070888
				11'd983: d_out <= 32'b00000000000000010001001001010010; // d_in = 2.919922, d_out = 1.071557
				11'd984: d_out <= 32'b00000000000000010001001001111101; // d_in = 2.921875, d_out = 1.072226
				11'd985: d_out <= 32'b00000000000000010001001010101001; // d_in = 2.923828, d_out = 1.072894
				11'd986: d_out <= 32'b00000000000000010001001011010101; // d_in = 2.925781, d_out = 1.073562
				11'd987: d_out <= 32'b00000000000000010001001100000001; // d_in = 2.927734, d_out = 1.074229
				11'd988: d_out <= 32'b00000000000000010001001100101100; // d_in = 2.929688, d_out = 1.074896
				11'd989: d_out <= 32'b00000000000000010001001101011000; // d_in = 2.931641, d_out = 1.075562
				11'd990: d_out <= 32'b00000000000000010001001110000100; // d_in = 2.933594, d_out = 1.076228
				11'd991: d_out <= 32'b00000000000000010001001110101111; // d_in = 2.935547, d_out = 1.076894
				11'd992: d_out <= 32'b00000000000000010001001111011011; // d_in = 2.937500, d_out = 1.077559
				11'd993: d_out <= 32'b00000000000000010001010000000110; // d_in = 2.939453, d_out = 1.078224
				11'd994: d_out <= 32'b00000000000000010001010000110010; // d_in = 2.941406, d_out = 1.078888
				11'd995: d_out <= 32'b00000000000000010001010001011101; // d_in = 2.943359, d_out = 1.079552
				11'd996: d_out <= 32'b00000000000000010001010010001001; // d_in = 2.945312, d_out = 1.080215
				11'd997: d_out <= 32'b00000000000000010001010010110100; // d_in = 2.947266, d_out = 1.080878
				11'd998: d_out <= 32'b00000000000000010001010011100000; // d_in = 2.949219, d_out = 1.081540
				11'd999: d_out <= 32'b00000000000000010001010100001011; // d_in = 2.951172, d_out = 1.082202
				11'd1000: d_out <= 32'b00000000000000010001010100110111; // d_in = 2.953125, d_out = 1.082864
				11'd1001: d_out <= 32'b00000000000000010001010101100010; // d_in = 2.955078, d_out = 1.083525
				11'd1002: d_out <= 32'b00000000000000010001010110001101; // d_in = 2.957031, d_out = 1.084186
				11'd1003: d_out <= 32'b00000000000000010001010110111000; // d_in = 2.958984, d_out = 1.084846
				11'd1004: d_out <= 32'b00000000000000010001010111100100; // d_in = 2.960938, d_out = 1.085506
				11'd1005: d_out <= 32'b00000000000000010001011000001111; // d_in = 2.962891, d_out = 1.086165
				11'd1006: d_out <= 32'b00000000000000010001011000111010; // d_in = 2.964844, d_out = 1.086824
				11'd1007: d_out <= 32'b00000000000000010001011001100101; // d_in = 2.966797, d_out = 1.087483
				11'd1008: d_out <= 32'b00000000000000010001011010010000; // d_in = 2.968750, d_out = 1.088141
				11'd1009: d_out <= 32'b00000000000000010001011010111100; // d_in = 2.970703, d_out = 1.088799
				11'd1010: d_out <= 32'b00000000000000010001011011100111; // d_in = 2.972656, d_out = 1.089456
				11'd1011: d_out <= 32'b00000000000000010001011100010010; // d_in = 2.974609, d_out = 1.090113
				11'd1012: d_out <= 32'b00000000000000010001011100111101; // d_in = 2.976562, d_out = 1.090769
				11'd1013: d_out <= 32'b00000000000000010001011101101000; // d_in = 2.978516, d_out = 1.091425
				11'd1014: d_out <= 32'b00000000000000010001011110010011; // d_in = 2.980469, d_out = 1.092081
				11'd1015: d_out <= 32'b00000000000000010001011110111110; // d_in = 2.982422, d_out = 1.092736
				11'd1016: d_out <= 32'b00000000000000010001011111101000; // d_in = 2.984375, d_out = 1.093390
				11'd1017: d_out <= 32'b00000000000000010001100000010011; // d_in = 2.986328, d_out = 1.094045
				11'd1018: d_out <= 32'b00000000000000010001100000111110; // d_in = 2.988281, d_out = 1.094698
				11'd1019: d_out <= 32'b00000000000000010001100001101001; // d_in = 2.990234, d_out = 1.095352
				11'd1020: d_out <= 32'b00000000000000010001100010010100; // d_in = 2.992188, d_out = 1.096005
				11'd1021: d_out <= 32'b00000000000000010001100010111111; // d_in = 2.994141, d_out = 1.096657
				11'd1022: d_out <= 32'b00000000000000010001100011101001; // d_in = 2.996094, d_out = 1.097309
				11'd1023: d_out <= 32'b00000000000000010001100100010100; // d_in = 2.998047, d_out = 1.097961
				11'd1024: d_out <= 32'b00000000000000010001100100111111; // d_in = 3.000000, d_out = 1.098612
				11'd1025: d_out <= 32'b00000000000000010001100101101001; // d_in = 3.001953, d_out = 1.099263
				11'd1026: d_out <= 32'b00000000000000010001100110010100; // d_in = 3.003906, d_out = 1.099914
				11'd1027: d_out <= 32'b00000000000000010001100110111111; // d_in = 3.005859, d_out = 1.100564
				11'd1028: d_out <= 32'b00000000000000010001100111101001; // d_in = 3.007812, d_out = 1.101213
				11'd1029: d_out <= 32'b00000000000000010001101000010100; // d_in = 3.009766, d_out = 1.101862
				11'd1030: d_out <= 32'b00000000000000010001101000111110; // d_in = 3.011719, d_out = 1.102511
				11'd1031: d_out <= 32'b00000000000000010001101001101001; // d_in = 3.013672, d_out = 1.103159
				11'd1032: d_out <= 32'b00000000000000010001101010010011; // d_in = 3.015625, d_out = 1.103807
				11'd1033: d_out <= 32'b00000000000000010001101010111110; // d_in = 3.017578, d_out = 1.104455
				11'd1034: d_out <= 32'b00000000000000010001101011101000; // d_in = 3.019531, d_out = 1.105102
				11'd1035: d_out <= 32'b00000000000000010001101100010010; // d_in = 3.021484, d_out = 1.105748
				11'd1036: d_out <= 32'b00000000000000010001101100111101; // d_in = 3.023438, d_out = 1.106394
				11'd1037: d_out <= 32'b00000000000000010001101101100111; // d_in = 3.025391, d_out = 1.107040
				11'd1038: d_out <= 32'b00000000000000010001101110010001; // d_in = 3.027344, d_out = 1.107686
				11'd1039: d_out <= 32'b00000000000000010001101110111100; // d_in = 3.029297, d_out = 1.108331
				11'd1040: d_out <= 32'b00000000000000010001101111100110; // d_in = 3.031250, d_out = 1.108975
				11'd1041: d_out <= 32'b00000000000000010001110000010000; // d_in = 3.033203, d_out = 1.109619
				11'd1042: d_out <= 32'b00000000000000010001110000111010; // d_in = 3.035156, d_out = 1.110263
				11'd1043: d_out <= 32'b00000000000000010001110001100100; // d_in = 3.037109, d_out = 1.110906
				11'd1044: d_out <= 32'b00000000000000010001110010001110; // d_in = 3.039062, d_out = 1.111549
				11'd1045: d_out <= 32'b00000000000000010001110010111001; // d_in = 3.041016, d_out = 1.112192
				11'd1046: d_out <= 32'b00000000000000010001110011100011; // d_in = 3.042969, d_out = 1.112834
				11'd1047: d_out <= 32'b00000000000000010001110100001101; // d_in = 3.044922, d_out = 1.113475
				11'd1048: d_out <= 32'b00000000000000010001110100110111; // d_in = 3.046875, d_out = 1.114116
				11'd1049: d_out <= 32'b00000000000000010001110101100001; // d_in = 3.048828, d_out = 1.114757
				11'd1050: d_out <= 32'b00000000000000010001110110001011; // d_in = 3.050781, d_out = 1.115398
				11'd1051: d_out <= 32'b00000000000000010001110110110101; // d_in = 3.052734, d_out = 1.116038
				11'd1052: d_out <= 32'b00000000000000010001110111011111; // d_in = 3.054688, d_out = 1.116677
				11'd1053: d_out <= 32'b00000000000000010001111000001000; // d_in = 3.056641, d_out = 1.117316
				11'd1054: d_out <= 32'b00000000000000010001111000110010; // d_in = 3.058594, d_out = 1.117955
				11'd1055: d_out <= 32'b00000000000000010001111001011100; // d_in = 3.060547, d_out = 1.118594
				11'd1056: d_out <= 32'b00000000000000010001111010000110; // d_in = 3.062500, d_out = 1.119232
				11'd1057: d_out <= 32'b00000000000000010001111010110000; // d_in = 3.064453, d_out = 1.119869
				11'd1058: d_out <= 32'b00000000000000010001111011011001; // d_in = 3.066406, d_out = 1.120506
				11'd1059: d_out <= 32'b00000000000000010001111100000011; // d_in = 3.068359, d_out = 1.121143
				11'd1060: d_out <= 32'b00000000000000010001111100101101; // d_in = 3.070312, d_out = 1.121779
				11'd1061: d_out <= 32'b00000000000000010001111101010111; // d_in = 3.072266, d_out = 1.122415
				11'd1062: d_out <= 32'b00000000000000010001111110000000; // d_in = 3.074219, d_out = 1.123051
				11'd1063: d_out <= 32'b00000000000000010001111110101010; // d_in = 3.076172, d_out = 1.123686
				11'd1064: d_out <= 32'b00000000000000010001111111010011; // d_in = 3.078125, d_out = 1.124321
				11'd1065: d_out <= 32'b00000000000000010001111111111101; // d_in = 3.080078, d_out = 1.124955
				11'd1066: d_out <= 32'b00000000000000010010000000100111; // d_in = 3.082031, d_out = 1.125589
				11'd1067: d_out <= 32'b00000000000000010010000001010000; // d_in = 3.083984, d_out = 1.126222
				11'd1068: d_out <= 32'b00000000000000010010000001111010; // d_in = 3.085938, d_out = 1.126856
				11'd1069: d_out <= 32'b00000000000000010010000010100011; // d_in = 3.087891, d_out = 1.127488
				11'd1070: d_out <= 32'b00000000000000010010000011001101; // d_in = 3.089844, d_out = 1.128121
				11'd1071: d_out <= 32'b00000000000000010010000011110110; // d_in = 3.091797, d_out = 1.128752
				11'd1072: d_out <= 32'b00000000000000010010000100011111; // d_in = 3.093750, d_out = 1.129384
				11'd1073: d_out <= 32'b00000000000000010010000101001001; // d_in = 3.095703, d_out = 1.130015
				11'd1074: d_out <= 32'b00000000000000010010000101110010; // d_in = 3.097656, d_out = 1.130646
				11'd1075: d_out <= 32'b00000000000000010010000110011011; // d_in = 3.099609, d_out = 1.131276
				11'd1076: d_out <= 32'b00000000000000010010000111000101; // d_in = 3.101562, d_out = 1.131906
				11'd1077: d_out <= 32'b00000000000000010010000111101110; // d_in = 3.103516, d_out = 1.132536
				11'd1078: d_out <= 32'b00000000000000010010001000010111; // d_in = 3.105469, d_out = 1.133165
				11'd1079: d_out <= 32'b00000000000000010010001001000000; // d_in = 3.107422, d_out = 1.133793
				11'd1080: d_out <= 32'b00000000000000010010001001101001; // d_in = 3.109375, d_out = 1.134422
				11'd1081: d_out <= 32'b00000000000000010010001010010011; // d_in = 3.111328, d_out = 1.135050
				11'd1082: d_out <= 32'b00000000000000010010001010111100; // d_in = 3.113281, d_out = 1.135677
				11'd1083: d_out <= 32'b00000000000000010010001011100101; // d_in = 3.115234, d_out = 1.136304
				11'd1084: d_out <= 32'b00000000000000010010001100001110; // d_in = 3.117188, d_out = 1.136931
				11'd1085: d_out <= 32'b00000000000000010010001100110111; // d_in = 3.119141, d_out = 1.137558
				11'd1086: d_out <= 32'b00000000000000010010001101100000; // d_in = 3.121094, d_out = 1.138184
				11'd1087: d_out <= 32'b00000000000000010010001110001001; // d_in = 3.123047, d_out = 1.138809
				11'd1088: d_out <= 32'b00000000000000010010001110110010; // d_in = 3.125000, d_out = 1.139434
				11'd1089: d_out <= 32'b00000000000000010010001111011011; // d_in = 3.126953, d_out = 1.140059
				11'd1090: d_out <= 32'b00000000000000010010010000000100; // d_in = 3.128906, d_out = 1.140684
				11'd1091: d_out <= 32'b00000000000000010010010000101101; // d_in = 3.130859, d_out = 1.141308
				11'd1092: d_out <= 32'b00000000000000010010010001010110; // d_in = 3.132812, d_out = 1.141931
				11'd1093: d_out <= 32'b00000000000000010010010001111110; // d_in = 3.134766, d_out = 1.142554
				11'd1094: d_out <= 32'b00000000000000010010010010100111; // d_in = 3.136719, d_out = 1.143177
				11'd1095: d_out <= 32'b00000000000000010010010011010000; // d_in = 3.138672, d_out = 1.143800
				11'd1096: d_out <= 32'b00000000000000010010010011111001; // d_in = 3.140625, d_out = 1.144422
				11'd1097: d_out <= 32'b00000000000000010010010100100010; // d_in = 3.142578, d_out = 1.145044
				11'd1098: d_out <= 32'b00000000000000010010010101001010; // d_in = 3.144531, d_out = 1.145665
				11'd1099: d_out <= 32'b00000000000000010010010101110011; // d_in = 3.146484, d_out = 1.146286
				11'd1100: d_out <= 32'b00000000000000010010010110011100; // d_in = 3.148438, d_out = 1.146906
				11'd1101: d_out <= 32'b00000000000000010010010111000100; // d_in = 3.150391, d_out = 1.147526
				11'd1102: d_out <= 32'b00000000000000010010010111101101; // d_in = 3.152344, d_out = 1.148146
				11'd1103: d_out <= 32'b00000000000000010010011000010110; // d_in = 3.154297, d_out = 1.148766
				11'd1104: d_out <= 32'b00000000000000010010011000111110; // d_in = 3.156250, d_out = 1.149385
				11'd1105: d_out <= 32'b00000000000000010010011001100111; // d_in = 3.158203, d_out = 1.150003
				11'd1106: d_out <= 32'b00000000000000010010011010001111; // d_in = 3.160156, d_out = 1.150621
				11'd1107: d_out <= 32'b00000000000000010010011010111000; // d_in = 3.162109, d_out = 1.151239
				11'd1108: d_out <= 32'b00000000000000010010011011100000; // d_in = 3.164062, d_out = 1.151857
				11'd1109: d_out <= 32'b00000000000000010010011100001001; // d_in = 3.166016, d_out = 1.152474
				11'd1110: d_out <= 32'b00000000000000010010011100110001; // d_in = 3.167969, d_out = 1.153091
				11'd1111: d_out <= 32'b00000000000000010010011101011001; // d_in = 3.169922, d_out = 1.153707
				11'd1112: d_out <= 32'b00000000000000010010011110000010; // d_in = 3.171875, d_out = 1.154323
				11'd1113: d_out <= 32'b00000000000000010010011110101010; // d_in = 3.173828, d_out = 1.154938
				11'd1114: d_out <= 32'b00000000000000010010011111010010; // d_in = 3.175781, d_out = 1.155554
				11'd1115: d_out <= 32'b00000000000000010010011111111011; // d_in = 3.177734, d_out = 1.156168
				11'd1116: d_out <= 32'b00000000000000010010100000100011; // d_in = 3.179688, d_out = 1.156783
				11'd1117: d_out <= 32'b00000000000000010010100001001011; // d_in = 3.181641, d_out = 1.157397
				11'd1118: d_out <= 32'b00000000000000010010100001110011; // d_in = 3.183594, d_out = 1.158011
				11'd1119: d_out <= 32'b00000000000000010010100010011100; // d_in = 3.185547, d_out = 1.158624
				11'd1120: d_out <= 32'b00000000000000010010100011000100; // d_in = 3.187500, d_out = 1.159237
				11'd1121: d_out <= 32'b00000000000000010010100011101100; // d_in = 3.189453, d_out = 1.159849
				11'd1122: d_out <= 32'b00000000000000010010100100010100; // d_in = 3.191406, d_out = 1.160462
				11'd1123: d_out <= 32'b00000000000000010010100100111100; // d_in = 3.193359, d_out = 1.161073
				11'd1124: d_out <= 32'b00000000000000010010100101100100; // d_in = 3.195312, d_out = 1.161685
				11'd1125: d_out <= 32'b00000000000000010010100110001100; // d_in = 3.197266, d_out = 1.162296
				11'd1126: d_out <= 32'b00000000000000010010100110110100; // d_in = 3.199219, d_out = 1.162907
				11'd1127: d_out <= 32'b00000000000000010010100111011100; // d_in = 3.201172, d_out = 1.163517
				11'd1128: d_out <= 32'b00000000000000010010101000000100; // d_in = 3.203125, d_out = 1.164127
				11'd1129: d_out <= 32'b00000000000000010010101000101100; // d_in = 3.205078, d_out = 1.164736
				11'd1130: d_out <= 32'b00000000000000010010101001010100; // d_in = 3.207031, d_out = 1.165346
				11'd1131: d_out <= 32'b00000000000000010010101001111100; // d_in = 3.208984, d_out = 1.165954
				11'd1132: d_out <= 32'b00000000000000010010101010100100; // d_in = 3.210938, d_out = 1.166563
				11'd1133: d_out <= 32'b00000000000000010010101011001100; // d_in = 3.212891, d_out = 1.167171
				11'd1134: d_out <= 32'b00000000000000010010101011110100; // d_in = 3.214844, d_out = 1.167779
				11'd1135: d_out <= 32'b00000000000000010010101100011011; // d_in = 3.216797, d_out = 1.168386
				11'd1136: d_out <= 32'b00000000000000010010101101000011; // d_in = 3.218750, d_out = 1.168993
				11'd1137: d_out <= 32'b00000000000000010010101101101011; // d_in = 3.220703, d_out = 1.169600
				11'd1138: d_out <= 32'b00000000000000010010101110010011; // d_in = 3.222656, d_out = 1.170206
				11'd1139: d_out <= 32'b00000000000000010010101110111010; // d_in = 3.224609, d_out = 1.170812
				11'd1140: d_out <= 32'b00000000000000010010101111100010; // d_in = 3.226562, d_out = 1.171417
				11'd1141: d_out <= 32'b00000000000000010010110000001010; // d_in = 3.228516, d_out = 1.172022
				11'd1142: d_out <= 32'b00000000000000010010110000110001; // d_in = 3.230469, d_out = 1.172627
				11'd1143: d_out <= 32'b00000000000000010010110001011001; // d_in = 3.232422, d_out = 1.173232
				11'd1144: d_out <= 32'b00000000000000010010110010000000; // d_in = 3.234375, d_out = 1.173836
				11'd1145: d_out <= 32'b00000000000000010010110010101000; // d_in = 3.236328, d_out = 1.174439
				11'd1146: d_out <= 32'b00000000000000010010110011010000; // d_in = 3.238281, d_out = 1.175043
				11'd1147: d_out <= 32'b00000000000000010010110011110111; // d_in = 3.240234, d_out = 1.175646
				11'd1148: d_out <= 32'b00000000000000010010110100011111; // d_in = 3.242188, d_out = 1.176248
				11'd1149: d_out <= 32'b00000000000000010010110101000110; // d_in = 3.244141, d_out = 1.176850
				11'd1150: d_out <= 32'b00000000000000010010110101101110; // d_in = 3.246094, d_out = 1.177452
				11'd1151: d_out <= 32'b00000000000000010010110110010101; // d_in = 3.248047, d_out = 1.178054
				11'd1152: d_out <= 32'b00000000000000010010110110111100; // d_in = 3.250000, d_out = 1.178655
				11'd1153: d_out <= 32'b00000000000000010010110111100100; // d_in = 3.251953, d_out = 1.179256
				11'd1154: d_out <= 32'b00000000000000010010111000001011; // d_in = 3.253906, d_out = 1.179856
				11'd1155: d_out <= 32'b00000000000000010010111000110010; // d_in = 3.255859, d_out = 1.180456
				11'd1156: d_out <= 32'b00000000000000010010111001011010; // d_in = 3.257812, d_out = 1.181056
				11'd1157: d_out <= 32'b00000000000000010010111010000001; // d_in = 3.259766, d_out = 1.181655
				11'd1158: d_out <= 32'b00000000000000010010111010101000; // d_in = 3.261719, d_out = 1.182254
				11'd1159: d_out <= 32'b00000000000000010010111011001111; // d_in = 3.263672, d_out = 1.182853
				11'd1160: d_out <= 32'b00000000000000010010111011110111; // d_in = 3.265625, d_out = 1.183451
				11'd1161: d_out <= 32'b00000000000000010010111100011110; // d_in = 3.267578, d_out = 1.184049
				11'd1162: d_out <= 32'b00000000000000010010111101000101; // d_in = 3.269531, d_out = 1.184647
				11'd1163: d_out <= 32'b00000000000000010010111101101100; // d_in = 3.271484, d_out = 1.185244
				11'd1164: d_out <= 32'b00000000000000010010111110010011; // d_in = 3.273438, d_out = 1.185841
				11'd1165: d_out <= 32'b00000000000000010010111110111010; // d_in = 3.275391, d_out = 1.186437
				11'd1166: d_out <= 32'b00000000000000010010111111100001; // d_in = 3.277344, d_out = 1.187033
				11'd1167: d_out <= 32'b00000000000000010011000000001000; // d_in = 3.279297, d_out = 1.187629
				11'd1168: d_out <= 32'b00000000000000010011000000101111; // d_in = 3.281250, d_out = 1.188224
				11'd1169: d_out <= 32'b00000000000000010011000001010110; // d_in = 3.283203, d_out = 1.188820
				11'd1170: d_out <= 32'b00000000000000010011000001111101; // d_in = 3.285156, d_out = 1.189414
				11'd1171: d_out <= 32'b00000000000000010011000010100100; // d_in = 3.287109, d_out = 1.190009
				11'd1172: d_out <= 32'b00000000000000010011000011001011; // d_in = 3.289062, d_out = 1.190603
				11'd1173: d_out <= 32'b00000000000000010011000011110010; // d_in = 3.291016, d_out = 1.191196
				11'd1174: d_out <= 32'b00000000000000010011000100011001; // d_in = 3.292969, d_out = 1.191790
				11'd1175: d_out <= 32'b00000000000000010011000101000000; // d_in = 3.294922, d_out = 1.192382
				11'd1176: d_out <= 32'b00000000000000010011000101100111; // d_in = 3.296875, d_out = 1.192975
				11'd1177: d_out <= 32'b00000000000000010011000110001110; // d_in = 3.298828, d_out = 1.193567
				11'd1178: d_out <= 32'b00000000000000010011000110110100; // d_in = 3.300781, d_out = 1.194159
				11'd1179: d_out <= 32'b00000000000000010011000111011011; // d_in = 3.302734, d_out = 1.194751
				11'd1180: d_out <= 32'b00000000000000010011001000000010; // d_in = 3.304688, d_out = 1.195342
				11'd1181: d_out <= 32'b00000000000000010011001000101001; // d_in = 3.306641, d_out = 1.195933
				11'd1182: d_out <= 32'b00000000000000010011001001001111; // d_in = 3.308594, d_out = 1.196523
				11'd1183: d_out <= 32'b00000000000000010011001001110110; // d_in = 3.310547, d_out = 1.197113
				11'd1184: d_out <= 32'b00000000000000010011001010011101; // d_in = 3.312500, d_out = 1.197703
				11'd1185: d_out <= 32'b00000000000000010011001011000011; // d_in = 3.314453, d_out = 1.198293
				11'd1186: d_out <= 32'b00000000000000010011001011101010; // d_in = 3.316406, d_out = 1.198882
				11'd1187: d_out <= 32'b00000000000000010011001100010000; // d_in = 3.318359, d_out = 1.199470
				11'd1188: d_out <= 32'b00000000000000010011001100110111; // d_in = 3.320312, d_out = 1.200059
				11'd1189: d_out <= 32'b00000000000000010011001101011110; // d_in = 3.322266, d_out = 1.200647
				11'd1190: d_out <= 32'b00000000000000010011001110000100; // d_in = 3.324219, d_out = 1.201235
				11'd1191: d_out <= 32'b00000000000000010011001110101011; // d_in = 3.326172, d_out = 1.201822
				11'd1192: d_out <= 32'b00000000000000010011001111010001; // d_in = 3.328125, d_out = 1.202409
				11'd1193: d_out <= 32'b00000000000000010011001111111000; // d_in = 3.330078, d_out = 1.202996
				11'd1194: d_out <= 32'b00000000000000010011010000011110; // d_in = 3.332031, d_out = 1.203582
				11'd1195: d_out <= 32'b00000000000000010011010001000100; // d_in = 3.333984, d_out = 1.204168
				11'd1196: d_out <= 32'b00000000000000010011010001101011; // d_in = 3.335938, d_out = 1.204754
				11'd1197: d_out <= 32'b00000000000000010011010010010001; // d_in = 3.337891, d_out = 1.205339
				11'd1198: d_out <= 32'b00000000000000010011010010110111; // d_in = 3.339844, d_out = 1.205924
				11'd1199: d_out <= 32'b00000000000000010011010011011110; // d_in = 3.341797, d_out = 1.206509
				11'd1200: d_out <= 32'b00000000000000010011010100000100; // d_in = 3.343750, d_out = 1.207093
				11'd1201: d_out <= 32'b00000000000000010011010100101010; // d_in = 3.345703, d_out = 1.207677
				11'd1202: d_out <= 32'b00000000000000010011010101010001; // d_in = 3.347656, d_out = 1.208260
				11'd1203: d_out <= 32'b00000000000000010011010101110111; // d_in = 3.349609, d_out = 1.208844
				11'd1204: d_out <= 32'b00000000000000010011010110011101; // d_in = 3.351562, d_out = 1.209427
				11'd1205: d_out <= 32'b00000000000000010011010111000011; // d_in = 3.353516, d_out = 1.210009
				11'd1206: d_out <= 32'b00000000000000010011010111101001; // d_in = 3.355469, d_out = 1.210591
				11'd1207: d_out <= 32'b00000000000000010011011000001111; // d_in = 3.357422, d_out = 1.211173
				11'd1208: d_out <= 32'b00000000000000010011011000110110; // d_in = 3.359375, d_out = 1.211755
				11'd1209: d_out <= 32'b00000000000000010011011001011100; // d_in = 3.361328, d_out = 1.212336
				11'd1210: d_out <= 32'b00000000000000010011011010000010; // d_in = 3.363281, d_out = 1.212917
				11'd1211: d_out <= 32'b00000000000000010011011010101000; // d_in = 3.365234, d_out = 1.213498
				11'd1212: d_out <= 32'b00000000000000010011011011001110; // d_in = 3.367188, d_out = 1.214078
				11'd1213: d_out <= 32'b00000000000000010011011011110100; // d_in = 3.369141, d_out = 1.214658
				11'd1214: d_out <= 32'b00000000000000010011011100011010; // d_in = 3.371094, d_out = 1.215237
				11'd1215: d_out <= 32'b00000000000000010011011101000000; // d_in = 3.373047, d_out = 1.215816
				11'd1216: d_out <= 32'b00000000000000010011011101100110; // d_in = 3.375000, d_out = 1.216395
				11'd1217: d_out <= 32'b00000000000000010011011110001100; // d_in = 3.376953, d_out = 1.216974
				11'd1218: d_out <= 32'b00000000000000010011011110110001; // d_in = 3.378906, d_out = 1.217552
				11'd1219: d_out <= 32'b00000000000000010011011111010111; // d_in = 3.380859, d_out = 1.218130
				11'd1220: d_out <= 32'b00000000000000010011011111111101; // d_in = 3.382812, d_out = 1.218707
				11'd1221: d_out <= 32'b00000000000000010011100000100011; // d_in = 3.384766, d_out = 1.219285
				11'd1222: d_out <= 32'b00000000000000010011100001001001; // d_in = 3.386719, d_out = 1.219862
				11'd1223: d_out <= 32'b00000000000000010011100001101111; // d_in = 3.388672, d_out = 1.220438
				11'd1224: d_out <= 32'b00000000000000010011100010010100; // d_in = 3.390625, d_out = 1.221014
				11'd1225: d_out <= 32'b00000000000000010011100010111010; // d_in = 3.392578, d_out = 1.221590
				11'd1226: d_out <= 32'b00000000000000010011100011100000; // d_in = 3.394531, d_out = 1.222166
				11'd1227: d_out <= 32'b00000000000000010011100100000110; // d_in = 3.396484, d_out = 1.222741
				11'd1228: d_out <= 32'b00000000000000010011100100101011; // d_in = 3.398438, d_out = 1.223316
				11'd1229: d_out <= 32'b00000000000000010011100101010001; // d_in = 3.400391, d_out = 1.223890
				11'd1230: d_out <= 32'b00000000000000010011100101110111; // d_in = 3.402344, d_out = 1.224465
				11'd1231: d_out <= 32'b00000000000000010011100110011100; // d_in = 3.404297, d_out = 1.225038
				11'd1232: d_out <= 32'b00000000000000010011100111000010; // d_in = 3.406250, d_out = 1.225612
				11'd1233: d_out <= 32'b00000000000000010011100111100111; // d_in = 3.408203, d_out = 1.226185
				11'd1234: d_out <= 32'b00000000000000010011101000001101; // d_in = 3.410156, d_out = 1.226758
				11'd1235: d_out <= 32'b00000000000000010011101000110010; // d_in = 3.412109, d_out = 1.227331
				11'd1236: d_out <= 32'b00000000000000010011101001011000; // d_in = 3.414062, d_out = 1.227903
				11'd1237: d_out <= 32'b00000000000000010011101001111101; // d_in = 3.416016, d_out = 1.228475
				11'd1238: d_out <= 32'b00000000000000010011101010100011; // d_in = 3.417969, d_out = 1.229046
				11'd1239: d_out <= 32'b00000000000000010011101011001000; // d_in = 3.419922, d_out = 1.229618
				11'd1240: d_out <= 32'b00000000000000010011101011101110; // d_in = 3.421875, d_out = 1.230189
				11'd1241: d_out <= 32'b00000000000000010011101100010011; // d_in = 3.423828, d_out = 1.230759
				11'd1242: d_out <= 32'b00000000000000010011101100111000; // d_in = 3.425781, d_out = 1.231330
				11'd1243: d_out <= 32'b00000000000000010011101101011110; // d_in = 3.427734, d_out = 1.231900
				11'd1244: d_out <= 32'b00000000000000010011101110000011; // d_in = 3.429688, d_out = 1.232469
				11'd1245: d_out <= 32'b00000000000000010011101110101000; // d_in = 3.431641, d_out = 1.233038
				11'd1246: d_out <= 32'b00000000000000010011101111001110; // d_in = 3.433594, d_out = 1.233607
				11'd1247: d_out <= 32'b00000000000000010011101111110011; // d_in = 3.435547, d_out = 1.234176
				11'd1248: d_out <= 32'b00000000000000010011110000011000; // d_in = 3.437500, d_out = 1.234744
				11'd1249: d_out <= 32'b00000000000000010011110000111101; // d_in = 3.439453, d_out = 1.235312
				11'd1250: d_out <= 32'b00000000000000010011110001100011; // d_in = 3.441406, d_out = 1.235880
				11'd1251: d_out <= 32'b00000000000000010011110010001000; // d_in = 3.443359, d_out = 1.236448
				11'd1252: d_out <= 32'b00000000000000010011110010101101; // d_in = 3.445312, d_out = 1.237015
				11'd1253: d_out <= 32'b00000000000000010011110011010010; // d_in = 3.447266, d_out = 1.237581
				11'd1254: d_out <= 32'b00000000000000010011110011110111; // d_in = 3.449219, d_out = 1.238148
				11'd1255: d_out <= 32'b00000000000000010011110100011100; // d_in = 3.451172, d_out = 1.238714
				11'd1256: d_out <= 32'b00000000000000010011110101000001; // d_in = 3.453125, d_out = 1.239280
				11'd1257: d_out <= 32'b00000000000000010011110101100110; // d_in = 3.455078, d_out = 1.239845
				11'd1258: d_out <= 32'b00000000000000010011110110001100; // d_in = 3.457031, d_out = 1.240410
				11'd1259: d_out <= 32'b00000000000000010011110110110001; // d_in = 3.458984, d_out = 1.240975
				11'd1260: d_out <= 32'b00000000000000010011110111010110; // d_in = 3.460938, d_out = 1.241540
				11'd1261: d_out <= 32'b00000000000000010011110111111011; // d_in = 3.462891, d_out = 1.242104
				11'd1262: d_out <= 32'b00000000000000010011111000011111; // d_in = 3.464844, d_out = 1.242668
				11'd1263: d_out <= 32'b00000000000000010011111001000100; // d_in = 3.466797, d_out = 1.243231
				11'd1264: d_out <= 32'b00000000000000010011111001101001; // d_in = 3.468750, d_out = 1.243794
				11'd1265: d_out <= 32'b00000000000000010011111010001110; // d_in = 3.470703, d_out = 1.244357
				11'd1266: d_out <= 32'b00000000000000010011111010110011; // d_in = 3.472656, d_out = 1.244920
				11'd1267: d_out <= 32'b00000000000000010011111011011000; // d_in = 3.474609, d_out = 1.245482
				11'd1268: d_out <= 32'b00000000000000010011111011111101; // d_in = 3.476562, d_out = 1.246044
				11'd1269: d_out <= 32'b00000000000000010011111100100010; // d_in = 3.478516, d_out = 1.246606
				11'd1270: d_out <= 32'b00000000000000010011111101000110; // d_in = 3.480469, d_out = 1.247167
				11'd1271: d_out <= 32'b00000000000000010011111101101011; // d_in = 3.482422, d_out = 1.247728
				11'd1272: d_out <= 32'b00000000000000010011111110010000; // d_in = 3.484375, d_out = 1.248289
				11'd1273: d_out <= 32'b00000000000000010011111110110101; // d_in = 3.486328, d_out = 1.248849
				11'd1274: d_out <= 32'b00000000000000010011111111011001; // d_in = 3.488281, d_out = 1.249409
				11'd1275: d_out <= 32'b00000000000000010011111111111110; // d_in = 3.490234, d_out = 1.249969
				11'd1276: d_out <= 32'b00000000000000010100000000100011; // d_in = 3.492188, d_out = 1.250528
				11'd1277: d_out <= 32'b00000000000000010100000001000111; // d_in = 3.494141, d_out = 1.251087
				11'd1278: d_out <= 32'b00000000000000010100000001101100; // d_in = 3.496094, d_out = 1.251646
				11'd1279: d_out <= 32'b00000000000000010100000010010000; // d_in = 3.498047, d_out = 1.252205
				11'd1280: d_out <= 32'b00000000000000010100000010110101; // d_in = 3.500000, d_out = 1.252763
				11'd1281: d_out <= 32'b00000000000000010100000011011010; // d_in = 3.501953, d_out = 1.253321
				11'd1282: d_out <= 32'b00000000000000010100000011111110; // d_in = 3.503906, d_out = 1.253878
				11'd1283: d_out <= 32'b00000000000000010100000100100011; // d_in = 3.505859, d_out = 1.254436
				11'd1284: d_out <= 32'b00000000000000010100000101000111; // d_in = 3.507812, d_out = 1.254993
				11'd1285: d_out <= 32'b00000000000000010100000101101100; // d_in = 3.509766, d_out = 1.255549
				11'd1286: d_out <= 32'b00000000000000010100000110010000; // d_in = 3.511719, d_out = 1.256106
				11'd1287: d_out <= 32'b00000000000000010100000110110101; // d_in = 3.513672, d_out = 1.256662
				11'd1288: d_out <= 32'b00000000000000010100000111011001; // d_in = 3.515625, d_out = 1.257217
				11'd1289: d_out <= 32'b00000000000000010100000111111101; // d_in = 3.517578, d_out = 1.257773
				11'd1290: d_out <= 32'b00000000000000010100001000100010; // d_in = 3.519531, d_out = 1.258328
				11'd1291: d_out <= 32'b00000000000000010100001001000110; // d_in = 3.521484, d_out = 1.258883
				11'd1292: d_out <= 32'b00000000000000010100001001101010; // d_in = 3.523438, d_out = 1.259437
				11'd1293: d_out <= 32'b00000000000000010100001010001111; // d_in = 3.525391, d_out = 1.259991
				11'd1294: d_out <= 32'b00000000000000010100001010110011; // d_in = 3.527344, d_out = 1.260545
				11'd1295: d_out <= 32'b00000000000000010100001011010111; // d_in = 3.529297, d_out = 1.261099
				11'd1296: d_out <= 32'b00000000000000010100001011111100; // d_in = 3.531250, d_out = 1.261652
				11'd1297: d_out <= 32'b00000000000000010100001100100000; // d_in = 3.533203, d_out = 1.262205
				11'd1298: d_out <= 32'b00000000000000010100001101000100; // d_in = 3.535156, d_out = 1.262757
				11'd1299: d_out <= 32'b00000000000000010100001101101000; // d_in = 3.537109, d_out = 1.263310
				11'd1300: d_out <= 32'b00000000000000010100001110001100; // d_in = 3.539062, d_out = 1.263862
				11'd1301: d_out <= 32'b00000000000000010100001110110001; // d_in = 3.541016, d_out = 1.264414
				11'd1302: d_out <= 32'b00000000000000010100001111010101; // d_in = 3.542969, d_out = 1.264965
				11'd1303: d_out <= 32'b00000000000000010100001111111001; // d_in = 3.544922, d_out = 1.265516
				11'd1304: d_out <= 32'b00000000000000010100010000011101; // d_in = 3.546875, d_out = 1.266067
				11'd1305: d_out <= 32'b00000000000000010100010001000001; // d_in = 3.548828, d_out = 1.266617
				11'd1306: d_out <= 32'b00000000000000010100010001100101; // d_in = 3.550781, d_out = 1.267168
				11'd1307: d_out <= 32'b00000000000000010100010010001001; // d_in = 3.552734, d_out = 1.267718
				11'd1308: d_out <= 32'b00000000000000010100010010101101; // d_in = 3.554688, d_out = 1.268267
				11'd1309: d_out <= 32'b00000000000000010100010011010001; // d_in = 3.556641, d_out = 1.268816
				11'd1310: d_out <= 32'b00000000000000010100010011110101; // d_in = 3.558594, d_out = 1.269365
				11'd1311: d_out <= 32'b00000000000000010100010100011001; // d_in = 3.560547, d_out = 1.269914
				11'd1312: d_out <= 32'b00000000000000010100010100111101; // d_in = 3.562500, d_out = 1.270463
				11'd1313: d_out <= 32'b00000000000000010100010101100001; // d_in = 3.564453, d_out = 1.271011
				11'd1314: d_out <= 32'b00000000000000010100010110000101; // d_in = 3.566406, d_out = 1.271558
				11'd1315: d_out <= 32'b00000000000000010100010110101001; // d_in = 3.568359, d_out = 1.272106
				11'd1316: d_out <= 32'b00000000000000010100010111001101; // d_in = 3.570312, d_out = 1.272653
				11'd1317: d_out <= 32'b00000000000000010100010111110000; // d_in = 3.572266, d_out = 1.273200
				11'd1318: d_out <= 32'b00000000000000010100011000010100; // d_in = 3.574219, d_out = 1.273747
				11'd1319: d_out <= 32'b00000000000000010100011000111000; // d_in = 3.576172, d_out = 1.274293
				11'd1320: d_out <= 32'b00000000000000010100011001011100; // d_in = 3.578125, d_out = 1.274839
				11'd1321: d_out <= 32'b00000000000000010100011010000000; // d_in = 3.580078, d_out = 1.275385
				11'd1322: d_out <= 32'b00000000000000010100011010100011; // d_in = 3.582031, d_out = 1.275930
				11'd1323: d_out <= 32'b00000000000000010100011011000111; // d_in = 3.583984, d_out = 1.276475
				11'd1324: d_out <= 32'b00000000000000010100011011101011; // d_in = 3.585938, d_out = 1.277020
				11'd1325: d_out <= 32'b00000000000000010100011100001110; // d_in = 3.587891, d_out = 1.277564
				11'd1326: d_out <= 32'b00000000000000010100011100110010; // d_in = 3.589844, d_out = 1.278109
				11'd1327: d_out <= 32'b00000000000000010100011101010110; // d_in = 3.591797, d_out = 1.278653
				11'd1328: d_out <= 32'b00000000000000010100011101111001; // d_in = 3.593750, d_out = 1.279196
				11'd1329: d_out <= 32'b00000000000000010100011110011101; // d_in = 3.595703, d_out = 1.279740
				11'd1330: d_out <= 32'b00000000000000010100011111000001; // d_in = 3.597656, d_out = 1.280283
				11'd1331: d_out <= 32'b00000000000000010100011111100100; // d_in = 3.599609, d_out = 1.280825
				11'd1332: d_out <= 32'b00000000000000010100100000001000; // d_in = 3.601562, d_out = 1.281368
				11'd1333: d_out <= 32'b00000000000000010100100000101011; // d_in = 3.603516, d_out = 1.281910
				11'd1334: d_out <= 32'b00000000000000010100100001001111; // d_in = 3.605469, d_out = 1.282452
				11'd1335: d_out <= 32'b00000000000000010100100001110010; // d_in = 3.607422, d_out = 1.282993
				11'd1336: d_out <= 32'b00000000000000010100100010010110; // d_in = 3.609375, d_out = 1.283535
				11'd1337: d_out <= 32'b00000000000000010100100010111001; // d_in = 3.611328, d_out = 1.284076
				11'd1338: d_out <= 32'b00000000000000010100100011011101; // d_in = 3.613281, d_out = 1.284616
				11'd1339: d_out <= 32'b00000000000000010100100100000000; // d_in = 3.615234, d_out = 1.285157
				11'd1340: d_out <= 32'b00000000000000010100100100100011; // d_in = 3.617188, d_out = 1.285697
				11'd1341: d_out <= 32'b00000000000000010100100101000111; // d_in = 3.619141, d_out = 1.286237
				11'd1342: d_out <= 32'b00000000000000010100100101101010; // d_in = 3.621094, d_out = 1.286776
				11'd1343: d_out <= 32'b00000000000000010100100110001101; // d_in = 3.623047, d_out = 1.287315
				11'd1344: d_out <= 32'b00000000000000010100100110110001; // d_in = 3.625000, d_out = 1.287854
				11'd1345: d_out <= 32'b00000000000000010100100111010100; // d_in = 3.626953, d_out = 1.288393
				11'd1346: d_out <= 32'b00000000000000010100100111110111; // d_in = 3.628906, d_out = 1.288931
				11'd1347: d_out <= 32'b00000000000000010100101000011011; // d_in = 3.630859, d_out = 1.289469
				11'd1348: d_out <= 32'b00000000000000010100101000111110; // d_in = 3.632812, d_out = 1.290007
				11'd1349: d_out <= 32'b00000000000000010100101001100001; // d_in = 3.634766, d_out = 1.290545
				11'd1350: d_out <= 32'b00000000000000010100101010000100; // d_in = 3.636719, d_out = 1.291082
				11'd1351: d_out <= 32'b00000000000000010100101010101000; // d_in = 3.638672, d_out = 1.291619
				11'd1352: d_out <= 32'b00000000000000010100101011001011; // d_in = 3.640625, d_out = 1.292155
				11'd1353: d_out <= 32'b00000000000000010100101011101110; // d_in = 3.642578, d_out = 1.292692
				11'd1354: d_out <= 32'b00000000000000010100101100010001; // d_in = 3.644531, d_out = 1.293228
				11'd1355: d_out <= 32'b00000000000000010100101100110100; // d_in = 3.646484, d_out = 1.293764
				11'd1356: d_out <= 32'b00000000000000010100101101010111; // d_in = 3.648438, d_out = 1.294299
				11'd1357: d_out <= 32'b00000000000000010100101101111010; // d_in = 3.650391, d_out = 1.294834
				11'd1358: d_out <= 32'b00000000000000010100101110011101; // d_in = 3.652344, d_out = 1.295369
				11'd1359: d_out <= 32'b00000000000000010100101111000000; // d_in = 3.654297, d_out = 1.295904
				11'd1360: d_out <= 32'b00000000000000010100101111100011; // d_in = 3.656250, d_out = 1.296438
				11'd1361: d_out <= 32'b00000000000000010100110000000110; // d_in = 3.658203, d_out = 1.296972
				11'd1362: d_out <= 32'b00000000000000010100110000101001; // d_in = 3.660156, d_out = 1.297506
				11'd1363: d_out <= 32'b00000000000000010100110001001100; // d_in = 3.662109, d_out = 1.298039
				11'd1364: d_out <= 32'b00000000000000010100110001101111; // d_in = 3.664062, d_out = 1.298573
				11'd1365: d_out <= 32'b00000000000000010100110010010010; // d_in = 3.666016, d_out = 1.299105
				11'd1366: d_out <= 32'b00000000000000010100110010110101; // d_in = 3.667969, d_out = 1.299638
				11'd1367: d_out <= 32'b00000000000000010100110011011000; // d_in = 3.669922, d_out = 1.300170
				11'd1368: d_out <= 32'b00000000000000010100110011111011; // d_in = 3.671875, d_out = 1.300702
				11'd1369: d_out <= 32'b00000000000000010100110100011110; // d_in = 3.673828, d_out = 1.301234
				11'd1370: d_out <= 32'b00000000000000010100110101000001; // d_in = 3.675781, d_out = 1.301766
				11'd1371: d_out <= 32'b00000000000000010100110101100011; // d_in = 3.677734, d_out = 1.302297
				11'd1372: d_out <= 32'b00000000000000010100110110000110; // d_in = 3.679688, d_out = 1.302828
				11'd1373: d_out <= 32'b00000000000000010100110110101001; // d_in = 3.681641, d_out = 1.303358
				11'd1374: d_out <= 32'b00000000000000010100110111001100; // d_in = 3.683594, d_out = 1.303889
				11'd1375: d_out <= 32'b00000000000000010100110111101110; // d_in = 3.685547, d_out = 1.304419
				11'd1376: d_out <= 32'b00000000000000010100111000010001; // d_in = 3.687500, d_out = 1.304949
				11'd1377: d_out <= 32'b00000000000000010100111000110100; // d_in = 3.689453, d_out = 1.305478
				11'd1378: d_out <= 32'b00000000000000010100111001010111; // d_in = 3.691406, d_out = 1.306007
				11'd1379: d_out <= 32'b00000000000000010100111001111001; // d_in = 3.693359, d_out = 1.306536
				11'd1380: d_out <= 32'b00000000000000010100111010011100; // d_in = 3.695312, d_out = 1.307065
				11'd1381: d_out <= 32'b00000000000000010100111010111110; // d_in = 3.697266, d_out = 1.307594
				11'd1382: d_out <= 32'b00000000000000010100111011100001; // d_in = 3.699219, d_out = 1.308122
				11'd1383: d_out <= 32'b00000000000000010100111100000100; // d_in = 3.701172, d_out = 1.308649
				11'd1384: d_out <= 32'b00000000000000010100111100100110; // d_in = 3.703125, d_out = 1.309177
				11'd1385: d_out <= 32'b00000000000000010100111101001001; // d_in = 3.705078, d_out = 1.309704
				11'd1386: d_out <= 32'b00000000000000010100111101101011; // d_in = 3.707031, d_out = 1.310231
				11'd1387: d_out <= 32'b00000000000000010100111110001110; // d_in = 3.708984, d_out = 1.310758
				11'd1388: d_out <= 32'b00000000000000010100111110110000; // d_in = 3.710938, d_out = 1.311285
				11'd1389: d_out <= 32'b00000000000000010100111111010011; // d_in = 3.712891, d_out = 1.311811
				11'd1390: d_out <= 32'b00000000000000010100111111110101; // d_in = 3.714844, d_out = 1.312337
				11'd1391: d_out <= 32'b00000000000000010101000000011000; // d_in = 3.716797, d_out = 1.312862
				11'd1392: d_out <= 32'b00000000000000010101000000111010; // d_in = 3.718750, d_out = 1.313388
				11'd1393: d_out <= 32'b00000000000000010101000001011101; // d_in = 3.720703, d_out = 1.313913
				11'd1394: d_out <= 32'b00000000000000010101000001111111; // d_in = 3.722656, d_out = 1.314437
				11'd1395: d_out <= 32'b00000000000000010101000010100001; // d_in = 3.724609, d_out = 1.314962
				11'd1396: d_out <= 32'b00000000000000010101000011000100; // d_in = 3.726562, d_out = 1.315486
				11'd1397: d_out <= 32'b00000000000000010101000011100110; // d_in = 3.728516, d_out = 1.316010
				11'd1398: d_out <= 32'b00000000000000010101000100001000; // d_in = 3.730469, d_out = 1.316534
				11'd1399: d_out <= 32'b00000000000000010101000100101011; // d_in = 3.732422, d_out = 1.317057
				11'd1400: d_out <= 32'b00000000000000010101000101001101; // d_in = 3.734375, d_out = 1.317580
				11'd1401: d_out <= 32'b00000000000000010101000101101111; // d_in = 3.736328, d_out = 1.318103
				11'd1402: d_out <= 32'b00000000000000010101000110010001; // d_in = 3.738281, d_out = 1.318626
				11'd1403: d_out <= 32'b00000000000000010101000110110100; // d_in = 3.740234, d_out = 1.319148
				11'd1404: d_out <= 32'b00000000000000010101000111010110; // d_in = 3.742188, d_out = 1.319670
				11'd1405: d_out <= 32'b00000000000000010101000111111000; // d_in = 3.744141, d_out = 1.320192
				11'd1406: d_out <= 32'b00000000000000010101001000011010; // d_in = 3.746094, d_out = 1.320714
				11'd1407: d_out <= 32'b00000000000000010101001000111100; // d_in = 3.748047, d_out = 1.321235
				11'd1408: d_out <= 32'b00000000000000010101001001011111; // d_in = 3.750000, d_out = 1.321756
				11'd1409: d_out <= 32'b00000000000000010101001010000001; // d_in = 3.751953, d_out = 1.322277
				11'd1410: d_out <= 32'b00000000000000010101001010100011; // d_in = 3.753906, d_out = 1.322797
				11'd1411: d_out <= 32'b00000000000000010101001011000101; // d_in = 3.755859, d_out = 1.323317
				11'd1412: d_out <= 32'b00000000000000010101001011100111; // d_in = 3.757812, d_out = 1.323837
				11'd1413: d_out <= 32'b00000000000000010101001100001001; // d_in = 3.759766, d_out = 1.324357
				11'd1414: d_out <= 32'b00000000000000010101001100101011; // d_in = 3.761719, d_out = 1.324876
				11'd1415: d_out <= 32'b00000000000000010101001101001101; // d_in = 3.763672, d_out = 1.325395
				11'd1416: d_out <= 32'b00000000000000010101001101101111; // d_in = 3.765625, d_out = 1.325914
				11'd1417: d_out <= 32'b00000000000000010101001110010001; // d_in = 3.767578, d_out = 1.326432
				11'd1418: d_out <= 32'b00000000000000010101001110110011; // d_in = 3.769531, d_out = 1.326951
				11'd1419: d_out <= 32'b00000000000000010101001111010101; // d_in = 3.771484, d_out = 1.327469
				11'd1420: d_out <= 32'b00000000000000010101001111110111; // d_in = 3.773438, d_out = 1.327986
				11'd1421: d_out <= 32'b00000000000000010101010000011001; // d_in = 3.775391, d_out = 1.328504
				11'd1422: d_out <= 32'b00000000000000010101010000111011; // d_in = 3.777344, d_out = 1.329021
				11'd1423: d_out <= 32'b00000000000000010101010001011101; // d_in = 3.779297, d_out = 1.329538
				11'd1424: d_out <= 32'b00000000000000010101010001111110; // d_in = 3.781250, d_out = 1.330055
				11'd1425: d_out <= 32'b00000000000000010101010010100000; // d_in = 3.783203, d_out = 1.330571
				11'd1426: d_out <= 32'b00000000000000010101010011000010; // d_in = 3.785156, d_out = 1.331087
				11'd1427: d_out <= 32'b00000000000000010101010011100100; // d_in = 3.787109, d_out = 1.331603
				11'd1428: d_out <= 32'b00000000000000010101010100000110; // d_in = 3.789062, d_out = 1.332119
				11'd1429: d_out <= 32'b00000000000000010101010100100111; // d_in = 3.791016, d_out = 1.332634
				11'd1430: d_out <= 32'b00000000000000010101010101001001; // d_in = 3.792969, d_out = 1.333149
				11'd1431: d_out <= 32'b00000000000000010101010101101011; // d_in = 3.794922, d_out = 1.333664
				11'd1432: d_out <= 32'b00000000000000010101010110001101; // d_in = 3.796875, d_out = 1.334178
				11'd1433: d_out <= 32'b00000000000000010101010110101110; // d_in = 3.798828, d_out = 1.334693
				11'd1434: d_out <= 32'b00000000000000010101010111010000; // d_in = 3.800781, d_out = 1.335207
				11'd1435: d_out <= 32'b00000000000000010101010111110010; // d_in = 3.802734, d_out = 1.335720
				11'd1436: d_out <= 32'b00000000000000010101011000010011; // d_in = 3.804688, d_out = 1.336234
				11'd1437: d_out <= 32'b00000000000000010101011000110101; // d_in = 3.806641, d_out = 1.336747
				11'd1438: d_out <= 32'b00000000000000010101011001010111; // d_in = 3.808594, d_out = 1.337260
				11'd1439: d_out <= 32'b00000000000000010101011001111000; // d_in = 3.810547, d_out = 1.337773
				11'd1440: d_out <= 32'b00000000000000010101011010011010; // d_in = 3.812500, d_out = 1.338285
				11'd1441: d_out <= 32'b00000000000000010101011010111011; // d_in = 3.814453, d_out = 1.338797
				11'd1442: d_out <= 32'b00000000000000010101011011011101; // d_in = 3.816406, d_out = 1.339309
				11'd1443: d_out <= 32'b00000000000000010101011011111110; // d_in = 3.818359, d_out = 1.339821
				11'd1444: d_out <= 32'b00000000000000010101011100100000; // d_in = 3.820312, d_out = 1.340332
				11'd1445: d_out <= 32'b00000000000000010101011101000010; // d_in = 3.822266, d_out = 1.340843
				11'd1446: d_out <= 32'b00000000000000010101011101100011; // d_in = 3.824219, d_out = 1.341354
				11'd1447: d_out <= 32'b00000000000000010101011110000100; // d_in = 3.826172, d_out = 1.341865
				11'd1448: d_out <= 32'b00000000000000010101011110100110; // d_in = 3.828125, d_out = 1.342375
				11'd1449: d_out <= 32'b00000000000000010101011111000111; // d_in = 3.830078, d_out = 1.342885
				11'd1450: d_out <= 32'b00000000000000010101011111101001; // d_in = 3.832031, d_out = 1.343395
				11'd1451: d_out <= 32'b00000000000000010101100000001010; // d_in = 3.833984, d_out = 1.343905
				11'd1452: d_out <= 32'b00000000000000010101100000101100; // d_in = 3.835938, d_out = 1.344414
				11'd1453: d_out <= 32'b00000000000000010101100001001101; // d_in = 3.837891, d_out = 1.344923
				11'd1454: d_out <= 32'b00000000000000010101100001101110; // d_in = 3.839844, d_out = 1.345432
				11'd1455: d_out <= 32'b00000000000000010101100010010000; // d_in = 3.841797, d_out = 1.345940
				11'd1456: d_out <= 32'b00000000000000010101100010110001; // d_in = 3.843750, d_out = 1.346448
				11'd1457: d_out <= 32'b00000000000000010101100011010010; // d_in = 3.845703, d_out = 1.346956
				11'd1458: d_out <= 32'b00000000000000010101100011110011; // d_in = 3.847656, d_out = 1.347464
				11'd1459: d_out <= 32'b00000000000000010101100100010101; // d_in = 3.849609, d_out = 1.347972
				11'd1460: d_out <= 32'b00000000000000010101100100110110; // d_in = 3.851562, d_out = 1.348479
				11'd1461: d_out <= 32'b00000000000000010101100101010111; // d_in = 3.853516, d_out = 1.348986
				11'd1462: d_out <= 32'b00000000000000010101100101111000; // d_in = 3.855469, d_out = 1.349493
				11'd1463: d_out <= 32'b00000000000000010101100110011010; // d_in = 3.857422, d_out = 1.349999
				11'd1464: d_out <= 32'b00000000000000010101100110111011; // d_in = 3.859375, d_out = 1.350505
				11'd1465: d_out <= 32'b00000000000000010101100111011100; // d_in = 3.861328, d_out = 1.351011
				11'd1466: d_out <= 32'b00000000000000010101100111111101; // d_in = 3.863281, d_out = 1.351517
				11'd1467: d_out <= 32'b00000000000000010101101000011110; // d_in = 3.865234, d_out = 1.352022
				11'd1468: d_out <= 32'b00000000000000010101101000111111; // d_in = 3.867188, d_out = 1.352527
				11'd1469: d_out <= 32'b00000000000000010101101001100000; // d_in = 3.869141, d_out = 1.353032
				11'd1470: d_out <= 32'b00000000000000010101101010000001; // d_in = 3.871094, d_out = 1.353537
				11'd1471: d_out <= 32'b00000000000000010101101010100010; // d_in = 3.873047, d_out = 1.354042
				11'd1472: d_out <= 32'b00000000000000010101101011000100; // d_in = 3.875000, d_out = 1.354546
				11'd1473: d_out <= 32'b00000000000000010101101011100101; // d_in = 3.876953, d_out = 1.355050
				11'd1474: d_out <= 32'b00000000000000010101101100000110; // d_in = 3.878906, d_out = 1.355553
				11'd1475: d_out <= 32'b00000000000000010101101100100111; // d_in = 3.880859, d_out = 1.356057
				11'd1476: d_out <= 32'b00000000000000010101101101001000; // d_in = 3.882812, d_out = 1.356560
				11'd1477: d_out <= 32'b00000000000000010101101101101000; // d_in = 3.884766, d_out = 1.357063
				11'd1478: d_out <= 32'b00000000000000010101101110001001; // d_in = 3.886719, d_out = 1.357565
				11'd1479: d_out <= 32'b00000000000000010101101110101010; // d_in = 3.888672, d_out = 1.358068
				11'd1480: d_out <= 32'b00000000000000010101101111001011; // d_in = 3.890625, d_out = 1.358570
				11'd1481: d_out <= 32'b00000000000000010101101111101100; // d_in = 3.892578, d_out = 1.359072
				11'd1482: d_out <= 32'b00000000000000010101110000001101; // d_in = 3.894531, d_out = 1.359573
				11'd1483: d_out <= 32'b00000000000000010101110000101110; // d_in = 3.896484, d_out = 1.360075
				11'd1484: d_out <= 32'b00000000000000010101110001001111; // d_in = 3.898438, d_out = 1.360576
				11'd1485: d_out <= 32'b00000000000000010101110001110000; // d_in = 3.900391, d_out = 1.361077
				11'd1486: d_out <= 32'b00000000000000010101110010010000; // d_in = 3.902344, d_out = 1.361577
				11'd1487: d_out <= 32'b00000000000000010101110010110001; // d_in = 3.904297, d_out = 1.362078
				11'd1488: d_out <= 32'b00000000000000010101110011010010; // d_in = 3.906250, d_out = 1.362578
				11'd1489: d_out <= 32'b00000000000000010101110011110011; // d_in = 3.908203, d_out = 1.363078
				11'd1490: d_out <= 32'b00000000000000010101110100010011; // d_in = 3.910156, d_out = 1.363577
				11'd1491: d_out <= 32'b00000000000000010101110100110100; // d_in = 3.912109, d_out = 1.364077
				11'd1492: d_out <= 32'b00000000000000010101110101010101; // d_in = 3.914062, d_out = 1.364576
				11'd1493: d_out <= 32'b00000000000000010101110101110110; // d_in = 3.916016, d_out = 1.365075
				11'd1494: d_out <= 32'b00000000000000010101110110010110; // d_in = 3.917969, d_out = 1.365573
				11'd1495: d_out <= 32'b00000000000000010101110110110111; // d_in = 3.919922, d_out = 1.366072
				11'd1496: d_out <= 32'b00000000000000010101110111011000; // d_in = 3.921875, d_out = 1.366570
				11'd1497: d_out <= 32'b00000000000000010101110111111000; // d_in = 3.923828, d_out = 1.367068
				11'd1498: d_out <= 32'b00000000000000010101111000011001; // d_in = 3.925781, d_out = 1.367565
				11'd1499: d_out <= 32'b00000000000000010101111000111001; // d_in = 3.927734, d_out = 1.368063
				11'd1500: d_out <= 32'b00000000000000010101111001011010; // d_in = 3.929688, d_out = 1.368560
				11'd1501: d_out <= 32'b00000000000000010101111001111011; // d_in = 3.931641, d_out = 1.369057
				11'd1502: d_out <= 32'b00000000000000010101111010011011; // d_in = 3.933594, d_out = 1.369553
				11'd1503: d_out <= 32'b00000000000000010101111010111100; // d_in = 3.935547, d_out = 1.370050
				11'd1504: d_out <= 32'b00000000000000010101111011011100; // d_in = 3.937500, d_out = 1.370546
				11'd1505: d_out <= 32'b00000000000000010101111011111101; // d_in = 3.939453, d_out = 1.371042
				11'd1506: d_out <= 32'b00000000000000010101111100011101; // d_in = 3.941406, d_out = 1.371538
				11'd1507: d_out <= 32'b00000000000000010101111100111110; // d_in = 3.943359, d_out = 1.372033
				11'd1508: d_out <= 32'b00000000000000010101111101011110; // d_in = 3.945312, d_out = 1.372528
				11'd1509: d_out <= 32'b00000000000000010101111101111110; // d_in = 3.947266, d_out = 1.373023
				11'd1510: d_out <= 32'b00000000000000010101111110011111; // d_in = 3.949219, d_out = 1.373518
				11'd1511: d_out <= 32'b00000000000000010101111110111111; // d_in = 3.951172, d_out = 1.374012
				11'd1512: d_out <= 32'b00000000000000010101111111100000; // d_in = 3.953125, d_out = 1.374506
				11'd1513: d_out <= 32'b00000000000000010110000000000000; // d_in = 3.955078, d_out = 1.375000
				11'd1514: d_out <= 32'b00000000000000010110000000100000; // d_in = 3.957031, d_out = 1.375494
				11'd1515: d_out <= 32'b00000000000000010110000001000001; // d_in = 3.958984, d_out = 1.375988
				11'd1516: d_out <= 32'b00000000000000010110000001100001; // d_in = 3.960938, d_out = 1.376481
				11'd1517: d_out <= 32'b00000000000000010110000010000001; // d_in = 3.962891, d_out = 1.376974
				11'd1518: d_out <= 32'b00000000000000010110000010100010; // d_in = 3.964844, d_out = 1.377466
				11'd1519: d_out <= 32'b00000000000000010110000011000010; // d_in = 3.966797, d_out = 1.377959
				11'd1520: d_out <= 32'b00000000000000010110000011100010; // d_in = 3.968750, d_out = 1.378451
				11'd1521: d_out <= 32'b00000000000000010110000100000010; // d_in = 3.970703, d_out = 1.378943
				11'd1522: d_out <= 32'b00000000000000010110000100100011; // d_in = 3.972656, d_out = 1.379435
				11'd1523: d_out <= 32'b00000000000000010110000101000011; // d_in = 3.974609, d_out = 1.379926
				11'd1524: d_out <= 32'b00000000000000010110000101100011; // d_in = 3.976562, d_out = 1.380418
				11'd1525: d_out <= 32'b00000000000000010110000110000011; // d_in = 3.978516, d_out = 1.380909
				11'd1526: d_out <= 32'b00000000000000010110000110100011; // d_in = 3.980469, d_out = 1.381400
				11'd1527: d_out <= 32'b00000000000000010110000111000100; // d_in = 3.982422, d_out = 1.381890
				11'd1528: d_out <= 32'b00000000000000010110000111100100; // d_in = 3.984375, d_out = 1.382380
				11'd1529: d_out <= 32'b00000000000000010110001000000100; // d_in = 3.986328, d_out = 1.382871
				11'd1530: d_out <= 32'b00000000000000010110001000100100; // d_in = 3.988281, d_out = 1.383360
				11'd1531: d_out <= 32'b00000000000000010110001001000100; // d_in = 3.990234, d_out = 1.383850
				11'd1532: d_out <= 32'b00000000000000010110001001100100; // d_in = 3.992188, d_out = 1.384339
				11'd1533: d_out <= 32'b00000000000000010110001010000100; // d_in = 3.994141, d_out = 1.384828
				11'd1534: d_out <= 32'b00000000000000010110001010100100; // d_in = 3.996094, d_out = 1.385317
				11'd1535: d_out <= 32'b00000000000000010110001011000100; // d_in = 3.998047, d_out = 1.385806
				11'd1536: d_out <= 32'b00000000000000010110001011100100; // d_in = 4.000000, d_out = 1.386294
				11'd1537: d_out <= 32'b00000000000000010110001100000100; // d_in = 4.001953, d_out = 1.386783
				11'd1538: d_out <= 32'b00000000000000010110001100100100; // d_in = 4.003906, d_out = 1.387270
				11'd1539: d_out <= 32'b00000000000000010110001101000100; // d_in = 4.005859, d_out = 1.387758
				11'd1540: d_out <= 32'b00000000000000010110001101100100; // d_in = 4.007812, d_out = 1.388246
				11'd1541: d_out <= 32'b00000000000000010110001110000100; // d_in = 4.009766, d_out = 1.388733
				11'd1542: d_out <= 32'b00000000000000010110001110100100; // d_in = 4.011719, d_out = 1.389220
				11'd1543: d_out <= 32'b00000000000000010110001111000100; // d_in = 4.013672, d_out = 1.389707
				11'd1544: d_out <= 32'b00000000000000010110001111100100; // d_in = 4.015625, d_out = 1.390193
				11'd1545: d_out <= 32'b00000000000000010110010000000100; // d_in = 4.017578, d_out = 1.390679
				11'd1546: d_out <= 32'b00000000000000010110010000100011; // d_in = 4.019531, d_out = 1.391165
				11'd1547: d_out <= 32'b00000000000000010110010001000011; // d_in = 4.021484, d_out = 1.391651
				11'd1548: d_out <= 32'b00000000000000010110010001100011; // d_in = 4.023438, d_out = 1.392137
				11'd1549: d_out <= 32'b00000000000000010110010010000011; // d_in = 4.025391, d_out = 1.392622
				11'd1550: d_out <= 32'b00000000000000010110010010100011; // d_in = 4.027344, d_out = 1.393107
				11'd1551: d_out <= 32'b00000000000000010110010011000010; // d_in = 4.029297, d_out = 1.393592
				11'd1552: d_out <= 32'b00000000000000010110010011100010; // d_in = 4.031250, d_out = 1.394077
				11'd1553: d_out <= 32'b00000000000000010110010100000010; // d_in = 4.033203, d_out = 1.394561
				11'd1554: d_out <= 32'b00000000000000010110010100100010; // d_in = 4.035156, d_out = 1.395045
				11'd1555: d_out <= 32'b00000000000000010110010101000001; // d_in = 4.037109, d_out = 1.395529
				11'd1556: d_out <= 32'b00000000000000010110010101100001; // d_in = 4.039062, d_out = 1.396013
				11'd1557: d_out <= 32'b00000000000000010110010110000001; // d_in = 4.041016, d_out = 1.396496
				11'd1558: d_out <= 32'b00000000000000010110010110100000; // d_in = 4.042969, d_out = 1.396979
				11'd1559: d_out <= 32'b00000000000000010110010111000000; // d_in = 4.044922, d_out = 1.397462
				11'd1560: d_out <= 32'b00000000000000010110010111100000; // d_in = 4.046875, d_out = 1.397945
				11'd1561: d_out <= 32'b00000000000000010110010111111111; // d_in = 4.048828, d_out = 1.398427
				11'd1562: d_out <= 32'b00000000000000010110011000011111; // d_in = 4.050781, d_out = 1.398910
				11'd1563: d_out <= 32'b00000000000000010110011000111111; // d_in = 4.052734, d_out = 1.399392
				11'd1564: d_out <= 32'b00000000000000010110011001011110; // d_in = 4.054688, d_out = 1.399874
				11'd1565: d_out <= 32'b00000000000000010110011001111110; // d_in = 4.056641, d_out = 1.400355
				11'd1566: d_out <= 32'b00000000000000010110011010011101; // d_in = 4.058594, d_out = 1.400837
				11'd1567: d_out <= 32'b00000000000000010110011010111101; // d_in = 4.060547, d_out = 1.401318
				11'd1568: d_out <= 32'b00000000000000010110011011011100; // d_in = 4.062500, d_out = 1.401799
				11'd1569: d_out <= 32'b00000000000000010110011011111100; // d_in = 4.064453, d_out = 1.402279
				11'd1570: d_out <= 32'b00000000000000010110011100011011; // d_in = 4.066406, d_out = 1.402760
				11'd1571: d_out <= 32'b00000000000000010110011100111011; // d_in = 4.068359, d_out = 1.403240
				11'd1572: d_out <= 32'b00000000000000010110011101011010; // d_in = 4.070312, d_out = 1.403720
				11'd1573: d_out <= 32'b00000000000000010110011101111010; // d_in = 4.072266, d_out = 1.404200
				11'd1574: d_out <= 32'b00000000000000010110011110011001; // d_in = 4.074219, d_out = 1.404679
				11'd1575: d_out <= 32'b00000000000000010110011110111000; // d_in = 4.076172, d_out = 1.405158
				11'd1576: d_out <= 32'b00000000000000010110011111011000; // d_in = 4.078125, d_out = 1.405637
				11'd1577: d_out <= 32'b00000000000000010110011111110111; // d_in = 4.080078, d_out = 1.406116
				11'd1578: d_out <= 32'b00000000000000010110100000010111; // d_in = 4.082031, d_out = 1.406595
				11'd1579: d_out <= 32'b00000000000000010110100000110110; // d_in = 4.083984, d_out = 1.407073
				11'd1580: d_out <= 32'b00000000000000010110100001010101; // d_in = 4.085938, d_out = 1.407551
				11'd1581: d_out <= 32'b00000000000000010110100001110101; // d_in = 4.087891, d_out = 1.408029
				11'd1582: d_out <= 32'b00000000000000010110100010010100; // d_in = 4.089844, d_out = 1.408507
				11'd1583: d_out <= 32'b00000000000000010110100010110011; // d_in = 4.091797, d_out = 1.408984
				11'd1584: d_out <= 32'b00000000000000010110100011010010; // d_in = 4.093750, d_out = 1.409461
				11'd1585: d_out <= 32'b00000000000000010110100011110010; // d_in = 4.095703, d_out = 1.409938
				11'd1586: d_out <= 32'b00000000000000010110100100010001; // d_in = 4.097656, d_out = 1.410415
				11'd1587: d_out <= 32'b00000000000000010110100100110000; // d_in = 4.099609, d_out = 1.410892
				11'd1588: d_out <= 32'b00000000000000010110100101001111; // d_in = 4.101562, d_out = 1.411368
				11'd1589: d_out <= 32'b00000000000000010110100101101111; // d_in = 4.103516, d_out = 1.411844
				11'd1590: d_out <= 32'b00000000000000010110100110001110; // d_in = 4.105469, d_out = 1.412320
				11'd1591: d_out <= 32'b00000000000000010110100110101101; // d_in = 4.107422, d_out = 1.412796
				11'd1592: d_out <= 32'b00000000000000010110100111001100; // d_in = 4.109375, d_out = 1.413271
				11'd1593: d_out <= 32'b00000000000000010110100111101011; // d_in = 4.111328, d_out = 1.413746
				11'd1594: d_out <= 32'b00000000000000010110101000001010; // d_in = 4.113281, d_out = 1.414221
				11'd1595: d_out <= 32'b00000000000000010110101000101010; // d_in = 4.115234, d_out = 1.414696
				11'd1596: d_out <= 32'b00000000000000010110101001001001; // d_in = 4.117188, d_out = 1.415170
				11'd1597: d_out <= 32'b00000000000000010110101001101000; // d_in = 4.119141, d_out = 1.415645
				11'd1598: d_out <= 32'b00000000000000010110101010000111; // d_in = 4.121094, d_out = 1.416119
				11'd1599: d_out <= 32'b00000000000000010110101010100110; // d_in = 4.123047, d_out = 1.416592
				11'd1600: d_out <= 32'b00000000000000010110101011000101; // d_in = 4.125000, d_out = 1.417066
				11'd1601: d_out <= 32'b00000000000000010110101011100100; // d_in = 4.126953, d_out = 1.417539
				11'd1602: d_out <= 32'b00000000000000010110101100000011; // d_in = 4.128906, d_out = 1.418013
				11'd1603: d_out <= 32'b00000000000000010110101100100010; // d_in = 4.130859, d_out = 1.418485
				11'd1604: d_out <= 32'b00000000000000010110101101000001; // d_in = 4.132812, d_out = 1.418958
				11'd1605: d_out <= 32'b00000000000000010110101101100000; // d_in = 4.134766, d_out = 1.419431
				11'd1606: d_out <= 32'b00000000000000010110101101111111; // d_in = 4.136719, d_out = 1.419903
				11'd1607: d_out <= 32'b00000000000000010110101110011110; // d_in = 4.138672, d_out = 1.420375
				11'd1608: d_out <= 32'b00000000000000010110101110111101; // d_in = 4.140625, d_out = 1.420847
				11'd1609: d_out <= 32'b00000000000000010110101111011100; // d_in = 4.142578, d_out = 1.421318
				11'd1610: d_out <= 32'b00000000000000010110101111111010; // d_in = 4.144531, d_out = 1.421790
				11'd1611: d_out <= 32'b00000000000000010110110000011001; // d_in = 4.146484, d_out = 1.422261
				11'd1612: d_out <= 32'b00000000000000010110110000111000; // d_in = 4.148438, d_out = 1.422732
				11'd1613: d_out <= 32'b00000000000000010110110001010111; // d_in = 4.150391, d_out = 1.423202
				11'd1614: d_out <= 32'b00000000000000010110110001110110; // d_in = 4.152344, d_out = 1.423673
				11'd1615: d_out <= 32'b00000000000000010110110010010101; // d_in = 4.154297, d_out = 1.424143
				11'd1616: d_out <= 32'b00000000000000010110110010110011; // d_in = 4.156250, d_out = 1.424613
				11'd1617: d_out <= 32'b00000000000000010110110011010010; // d_in = 4.158203, d_out = 1.425083
				11'd1618: d_out <= 32'b00000000000000010110110011110001; // d_in = 4.160156, d_out = 1.425553
				11'd1619: d_out <= 32'b00000000000000010110110100010000; // d_in = 4.162109, d_out = 1.426022
				11'd1620: d_out <= 32'b00000000000000010110110100101111; // d_in = 4.164062, d_out = 1.426491
				11'd1621: d_out <= 32'b00000000000000010110110101001101; // d_in = 4.166016, d_out = 1.426960
				11'd1622: d_out <= 32'b00000000000000010110110101101100; // d_in = 4.167969, d_out = 1.427429
				11'd1623: d_out <= 32'b00000000000000010110110110001011; // d_in = 4.169922, d_out = 1.427897
				11'd1624: d_out <= 32'b00000000000000010110110110101001; // d_in = 4.171875, d_out = 1.428366
				11'd1625: d_out <= 32'b00000000000000010110110111001000; // d_in = 4.173828, d_out = 1.428834
				11'd1626: d_out <= 32'b00000000000000010110110111100111; // d_in = 4.175781, d_out = 1.429301
				11'd1627: d_out <= 32'b00000000000000010110111000000101; // d_in = 4.177734, d_out = 1.429769
				11'd1628: d_out <= 32'b00000000000000010110111000100100; // d_in = 4.179688, d_out = 1.430236
				11'd1629: d_out <= 32'b00000000000000010110111001000011; // d_in = 4.181641, d_out = 1.430704
				11'd1630: d_out <= 32'b00000000000000010110111001100001; // d_in = 4.183594, d_out = 1.431171
				11'd1631: d_out <= 32'b00000000000000010110111010000000; // d_in = 4.185547, d_out = 1.431637
				11'd1632: d_out <= 32'b00000000000000010110111010011110; // d_in = 4.187500, d_out = 1.432104
				11'd1633: d_out <= 32'b00000000000000010110111010111101; // d_in = 4.189453, d_out = 1.432570
				11'd1634: d_out <= 32'b00000000000000010110111011011011; // d_in = 4.191406, d_out = 1.433036
				11'd1635: d_out <= 32'b00000000000000010110111011111010; // d_in = 4.193359, d_out = 1.433502
				11'd1636: d_out <= 32'b00000000000000010110111100011001; // d_in = 4.195312, d_out = 1.433968
				11'd1637: d_out <= 32'b00000000000000010110111100110111; // d_in = 4.197266, d_out = 1.434433
				11'd1638: d_out <= 32'b00000000000000010110111101010110; // d_in = 4.199219, d_out = 1.434898
				11'd1639: d_out <= 32'b00000000000000010110111101110100; // d_in = 4.201172, d_out = 1.435364
				11'd1640: d_out <= 32'b00000000000000010110111110010010; // d_in = 4.203125, d_out = 1.435828
				11'd1641: d_out <= 32'b00000000000000010110111110110001; // d_in = 4.205078, d_out = 1.436293
				11'd1642: d_out <= 32'b00000000000000010110111111001111; // d_in = 4.207031, d_out = 1.436757
				11'd1643: d_out <= 32'b00000000000000010110111111101110; // d_in = 4.208984, d_out = 1.437221
				11'd1644: d_out <= 32'b00000000000000010111000000001100; // d_in = 4.210938, d_out = 1.437685
				11'd1645: d_out <= 32'b00000000000000010111000000101011; // d_in = 4.212891, d_out = 1.438149
				11'd1646: d_out <= 32'b00000000000000010111000001001001; // d_in = 4.214844, d_out = 1.438613
				11'd1647: d_out <= 32'b00000000000000010111000001100111; // d_in = 4.216797, d_out = 1.439076
				11'd1648: d_out <= 32'b00000000000000010111000010000110; // d_in = 4.218750, d_out = 1.439539
				11'd1649: d_out <= 32'b00000000000000010111000010100100; // d_in = 4.220703, d_out = 1.440002
				11'd1650: d_out <= 32'b00000000000000010111000011000010; // d_in = 4.222656, d_out = 1.440464
				11'd1651: d_out <= 32'b00000000000000010111000011100001; // d_in = 4.224609, d_out = 1.440927
				11'd1652: d_out <= 32'b00000000000000010111000011111111; // d_in = 4.226562, d_out = 1.441389
				11'd1653: d_out <= 32'b00000000000000010111000100011101; // d_in = 4.228516, d_out = 1.441851
				11'd1654: d_out <= 32'b00000000000000010111000100111011; // d_in = 4.230469, d_out = 1.442313
				11'd1655: d_out <= 32'b00000000000000010111000101011010; // d_in = 4.232422, d_out = 1.442774
				11'd1656: d_out <= 32'b00000000000000010111000101111000; // d_in = 4.234375, d_out = 1.443236
				11'd1657: d_out <= 32'b00000000000000010111000110010110; // d_in = 4.236328, d_out = 1.443697
				11'd1658: d_out <= 32'b00000000000000010111000110110100; // d_in = 4.238281, d_out = 1.444158
				11'd1659: d_out <= 32'b00000000000000010111000111010011; // d_in = 4.240234, d_out = 1.444619
				11'd1660: d_out <= 32'b00000000000000010111000111110001; // d_in = 4.242188, d_out = 1.445079
				11'd1661: d_out <= 32'b00000000000000010111001000001111; // d_in = 4.244141, d_out = 1.445539
				11'd1662: d_out <= 32'b00000000000000010111001000101101; // d_in = 4.246094, d_out = 1.445999
				11'd1663: d_out <= 32'b00000000000000010111001001001011; // d_in = 4.248047, d_out = 1.446459
				11'd1664: d_out <= 32'b00000000000000010111001001101001; // d_in = 4.250000, d_out = 1.446919
				11'd1665: d_out <= 32'b00000000000000010111001010000111; // d_in = 4.251953, d_out = 1.447378
				11'd1666: d_out <= 32'b00000000000000010111001010100101; // d_in = 4.253906, d_out = 1.447838
				11'd1667: d_out <= 32'b00000000000000010111001011000100; // d_in = 4.255859, d_out = 1.448297
				11'd1668: d_out <= 32'b00000000000000010111001011100010; // d_in = 4.257812, d_out = 1.448756
				11'd1669: d_out <= 32'b00000000000000010111001100000000; // d_in = 4.259766, d_out = 1.449214
				11'd1670: d_out <= 32'b00000000000000010111001100011110; // d_in = 4.261719, d_out = 1.449673
				11'd1671: d_out <= 32'b00000000000000010111001100111100; // d_in = 4.263672, d_out = 1.450131
				11'd1672: d_out <= 32'b00000000000000010111001101011010; // d_in = 4.265625, d_out = 1.450589
				11'd1673: d_out <= 32'b00000000000000010111001101111000; // d_in = 4.267578, d_out = 1.451046
				11'd1674: d_out <= 32'b00000000000000010111001110010110; // d_in = 4.269531, d_out = 1.451504
				11'd1675: d_out <= 32'b00000000000000010111001110110100; // d_in = 4.271484, d_out = 1.451961
				11'd1676: d_out <= 32'b00000000000000010111001111010010; // d_in = 4.273438, d_out = 1.452419
				11'd1677: d_out <= 32'b00000000000000010111001111110000; // d_in = 4.275391, d_out = 1.452875
				11'd1678: d_out <= 32'b00000000000000010111010000001110; // d_in = 4.277344, d_out = 1.453332
				11'd1679: d_out <= 32'b00000000000000010111010000101011; // d_in = 4.279297, d_out = 1.453789
				11'd1680: d_out <= 32'b00000000000000010111010001001001; // d_in = 4.281250, d_out = 1.454245
				11'd1681: d_out <= 32'b00000000000000010111010001100111; // d_in = 4.283203, d_out = 1.454701
				11'd1682: d_out <= 32'b00000000000000010111010010000101; // d_in = 4.285156, d_out = 1.455157
				11'd1683: d_out <= 32'b00000000000000010111010010100011; // d_in = 4.287109, d_out = 1.455613
				11'd1684: d_out <= 32'b00000000000000010111010011000001; // d_in = 4.289062, d_out = 1.456068
				11'd1685: d_out <= 32'b00000000000000010111010011011111; // d_in = 4.291016, d_out = 1.456523
				11'd1686: d_out <= 32'b00000000000000010111010011111101; // d_in = 4.292969, d_out = 1.456979
				11'd1687: d_out <= 32'b00000000000000010111010100011010; // d_in = 4.294922, d_out = 1.457433
				11'd1688: d_out <= 32'b00000000000000010111010100111000; // d_in = 4.296875, d_out = 1.457888
				11'd1689: d_out <= 32'b00000000000000010111010101010110; // d_in = 4.298828, d_out = 1.458342
				11'd1690: d_out <= 32'b00000000000000010111010101110100; // d_in = 4.300781, d_out = 1.458797
				11'd1691: d_out <= 32'b00000000000000010111010110010001; // d_in = 4.302734, d_out = 1.459251
				11'd1692: d_out <= 32'b00000000000000010111010110101111; // d_in = 4.304688, d_out = 1.459705
				11'd1693: d_out <= 32'b00000000000000010111010111001101; // d_in = 4.306641, d_out = 1.460158
				11'd1694: d_out <= 32'b00000000000000010111010111101011; // d_in = 4.308594, d_out = 1.460612
				11'd1695: d_out <= 32'b00000000000000010111011000001000; // d_in = 4.310547, d_out = 1.461065
				11'd1696: d_out <= 32'b00000000000000010111011000100110; // d_in = 4.312500, d_out = 1.461518
				11'd1697: d_out <= 32'b00000000000000010111011001000100; // d_in = 4.314453, d_out = 1.461971
				11'd1698: d_out <= 32'b00000000000000010111011001100001; // d_in = 4.316406, d_out = 1.462423
				11'd1699: d_out <= 32'b00000000000000010111011001111111; // d_in = 4.318359, d_out = 1.462876
				11'd1700: d_out <= 32'b00000000000000010111011010011101; // d_in = 4.320312, d_out = 1.463328
				11'd1701: d_out <= 32'b00000000000000010111011010111010; // d_in = 4.322266, d_out = 1.463780
				11'd1702: d_out <= 32'b00000000000000010111011011011000; // d_in = 4.324219, d_out = 1.464231
				11'd1703: d_out <= 32'b00000000000000010111011011110101; // d_in = 4.326172, d_out = 1.464683
				11'd1704: d_out <= 32'b00000000000000010111011100010011; // d_in = 4.328125, d_out = 1.465134
				11'd1705: d_out <= 32'b00000000000000010111011100110001; // d_in = 4.330078, d_out = 1.465586
				11'd1706: d_out <= 32'b00000000000000010111011101001110; // d_in = 4.332031, d_out = 1.466037
				11'd1707: d_out <= 32'b00000000000000010111011101101100; // d_in = 4.333984, d_out = 1.466487
				11'd1708: d_out <= 32'b00000000000000010111011110001001; // d_in = 4.335938, d_out = 1.466938
				11'd1709: d_out <= 32'b00000000000000010111011110100111; // d_in = 4.337891, d_out = 1.467388
				11'd1710: d_out <= 32'b00000000000000010111011111000100; // d_in = 4.339844, d_out = 1.467838
				11'd1711: d_out <= 32'b00000000000000010111011111100010; // d_in = 4.341797, d_out = 1.468288
				11'd1712: d_out <= 32'b00000000000000010111011111111111; // d_in = 4.343750, d_out = 1.468738
				11'd1713: d_out <= 32'b00000000000000010111100000011101; // d_in = 4.345703, d_out = 1.469188
				11'd1714: d_out <= 32'b00000000000000010111100000111010; // d_in = 4.347656, d_out = 1.469637
				11'd1715: d_out <= 32'b00000000000000010111100001011000; // d_in = 4.349609, d_out = 1.470086
				11'd1716: d_out <= 32'b00000000000000010111100001110101; // d_in = 4.351562, d_out = 1.470535
				11'd1717: d_out <= 32'b00000000000000010111100010010010; // d_in = 4.353516, d_out = 1.470984
				11'd1718: d_out <= 32'b00000000000000010111100010110000; // d_in = 4.355469, d_out = 1.471432
				11'd1719: d_out <= 32'b00000000000000010111100011001101; // d_in = 4.357422, d_out = 1.471881
				11'd1720: d_out <= 32'b00000000000000010111100011101011; // d_in = 4.359375, d_out = 1.472329
				11'd1721: d_out <= 32'b00000000000000010111100100001000; // d_in = 4.361328, d_out = 1.472777
				11'd1722: d_out <= 32'b00000000000000010111100100100101; // d_in = 4.363281, d_out = 1.473224
				11'd1723: d_out <= 32'b00000000000000010111100101000011; // d_in = 4.365234, d_out = 1.473672
				11'd1724: d_out <= 32'b00000000000000010111100101100000; // d_in = 4.367188, d_out = 1.474119
				11'd1725: d_out <= 32'b00000000000000010111100101111101; // d_in = 4.369141, d_out = 1.474566
				11'd1726: d_out <= 32'b00000000000000010111100110011010; // d_in = 4.371094, d_out = 1.475013
				11'd1727: d_out <= 32'b00000000000000010111100110111000; // d_in = 4.373047, d_out = 1.475460
				11'd1728: d_out <= 32'b00000000000000010111100111010101; // d_in = 4.375000, d_out = 1.475907
				11'd1729: d_out <= 32'b00000000000000010111100111110010; // d_in = 4.376953, d_out = 1.476353
				11'd1730: d_out <= 32'b00000000000000010111101000001111; // d_in = 4.378906, d_out = 1.476799
				11'd1731: d_out <= 32'b00000000000000010111101000101101; // d_in = 4.380859, d_out = 1.477245
				11'd1732: d_out <= 32'b00000000000000010111101001001010; // d_in = 4.382812, d_out = 1.477691
				11'd1733: d_out <= 32'b00000000000000010111101001100111; // d_in = 4.384766, d_out = 1.478136
				11'd1734: d_out <= 32'b00000000000000010111101010000100; // d_in = 4.386719, d_out = 1.478582
				11'd1735: d_out <= 32'b00000000000000010111101010100001; // d_in = 4.388672, d_out = 1.479027
				11'd1736: d_out <= 32'b00000000000000010111101010111111; // d_in = 4.390625, d_out = 1.479472
				11'd1737: d_out <= 32'b00000000000000010111101011011100; // d_in = 4.392578, d_out = 1.479916
				11'd1738: d_out <= 32'b00000000000000010111101011111001; // d_in = 4.394531, d_out = 1.480361
				11'd1739: d_out <= 32'b00000000000000010111101100010110; // d_in = 4.396484, d_out = 1.480805
				11'd1740: d_out <= 32'b00000000000000010111101100110011; // d_in = 4.398438, d_out = 1.481249
				11'd1741: d_out <= 32'b00000000000000010111101101010000; // d_in = 4.400391, d_out = 1.481693
				11'd1742: d_out <= 32'b00000000000000010111101101101101; // d_in = 4.402344, d_out = 1.482137
				11'd1743: d_out <= 32'b00000000000000010111101110001010; // d_in = 4.404297, d_out = 1.482581
				11'd1744: d_out <= 32'b00000000000000010111101110100111; // d_in = 4.406250, d_out = 1.483024
				11'd1745: d_out <= 32'b00000000000000010111101111000101; // d_in = 4.408203, d_out = 1.483467
				11'd1746: d_out <= 32'b00000000000000010111101111100010; // d_in = 4.410156, d_out = 1.483910
				11'd1747: d_out <= 32'b00000000000000010111101111111111; // d_in = 4.412109, d_out = 1.484353
				11'd1748: d_out <= 32'b00000000000000010111110000011100; // d_in = 4.414062, d_out = 1.484795
				11'd1749: d_out <= 32'b00000000000000010111110000111001; // d_in = 4.416016, d_out = 1.485238
				11'd1750: d_out <= 32'b00000000000000010111110001010110; // d_in = 4.417969, d_out = 1.485680
				11'd1751: d_out <= 32'b00000000000000010111110001110010; // d_in = 4.419922, d_out = 1.486122
				11'd1752: d_out <= 32'b00000000000000010111110010001111; // d_in = 4.421875, d_out = 1.486564
				11'd1753: d_out <= 32'b00000000000000010111110010101100; // d_in = 4.423828, d_out = 1.487005
				11'd1754: d_out <= 32'b00000000000000010111110011001001; // d_in = 4.425781, d_out = 1.487447
				11'd1755: d_out <= 32'b00000000000000010111110011100110; // d_in = 4.427734, d_out = 1.487888
				11'd1756: d_out <= 32'b00000000000000010111110100000011; // d_in = 4.429688, d_out = 1.488329
				11'd1757: d_out <= 32'b00000000000000010111110100100000; // d_in = 4.431641, d_out = 1.488770
				11'd1758: d_out <= 32'b00000000000000010111110100111101; // d_in = 4.433594, d_out = 1.489210
				11'd1759: d_out <= 32'b00000000000000010111110101011010; // d_in = 4.435547, d_out = 1.489651
				11'd1760: d_out <= 32'b00000000000000010111110101110111; // d_in = 4.437500, d_out = 1.490091
				11'd1761: d_out <= 32'b00000000000000010111110110010011; // d_in = 4.439453, d_out = 1.490531
				11'd1762: d_out <= 32'b00000000000000010111110110110000; // d_in = 4.441406, d_out = 1.490971
				11'd1763: d_out <= 32'b00000000000000010111110111001101; // d_in = 4.443359, d_out = 1.491411
				11'd1764: d_out <= 32'b00000000000000010111110111101010; // d_in = 4.445312, d_out = 1.491850
				11'd1765: d_out <= 32'b00000000000000010111111000000111; // d_in = 4.447266, d_out = 1.492289
				11'd1766: d_out <= 32'b00000000000000010111111000100011; // d_in = 4.449219, d_out = 1.492729
				11'd1767: d_out <= 32'b00000000000000010111111001000000; // d_in = 4.451172, d_out = 1.493167
				11'd1768: d_out <= 32'b00000000000000010111111001011101; // d_in = 4.453125, d_out = 1.493606
				11'd1769: d_out <= 32'b00000000000000010111111001111010; // d_in = 4.455078, d_out = 1.494045
				11'd1770: d_out <= 32'b00000000000000010111111010010110; // d_in = 4.457031, d_out = 1.494483
				11'd1771: d_out <= 32'b00000000000000010111111010110011; // d_in = 4.458984, d_out = 1.494921
				11'd1772: d_out <= 32'b00000000000000010111111011010000; // d_in = 4.460938, d_out = 1.495359
				11'd1773: d_out <= 32'b00000000000000010111111011101101; // d_in = 4.462891, d_out = 1.495797
				11'd1774: d_out <= 32'b00000000000000010111111100001001; // d_in = 4.464844, d_out = 1.496234
				11'd1775: d_out <= 32'b00000000000000010111111100100110; // d_in = 4.466797, d_out = 1.496672
				11'd1776: d_out <= 32'b00000000000000010111111101000011; // d_in = 4.468750, d_out = 1.497109
				11'd1777: d_out <= 32'b00000000000000010111111101011111; // d_in = 4.470703, d_out = 1.497546
				11'd1778: d_out <= 32'b00000000000000010111111101111100; // d_in = 4.472656, d_out = 1.497982
				11'd1779: d_out <= 32'b00000000000000010111111110011000; // d_in = 4.474609, d_out = 1.498419
				11'd1780: d_out <= 32'b00000000000000010111111110110101; // d_in = 4.476562, d_out = 1.498855
				11'd1781: d_out <= 32'b00000000000000010111111111010010; // d_in = 4.478516, d_out = 1.499292
				11'd1782: d_out <= 32'b00000000000000010111111111101110; // d_in = 4.480469, d_out = 1.499728
				11'd1783: d_out <= 32'b00000000000000011000000000001011; // d_in = 4.482422, d_out = 1.500163
				11'd1784: d_out <= 32'b00000000000000011000000000100111; // d_in = 4.484375, d_out = 1.500599
				11'd1785: d_out <= 32'b00000000000000011000000001000100; // d_in = 4.486328, d_out = 1.501035
				11'd1786: d_out <= 32'b00000000000000011000000001100000; // d_in = 4.488281, d_out = 1.501470
				11'd1787: d_out <= 32'b00000000000000011000000001111101; // d_in = 4.490234, d_out = 1.501905
				11'd1788: d_out <= 32'b00000000000000011000000010011001; // d_in = 4.492188, d_out = 1.502340
				11'd1789: d_out <= 32'b00000000000000011000000010110110; // d_in = 4.494141, d_out = 1.502774
				11'd1790: d_out <= 32'b00000000000000011000000011010010; // d_in = 4.496094, d_out = 1.503209
				11'd1791: d_out <= 32'b00000000000000011000000011101111; // d_in = 4.498047, d_out = 1.503643
				11'd1792: d_out <= 32'b00000000000000011000000100001011; // d_in = 4.500000, d_out = 1.504077
				11'd1793: d_out <= 32'b00000000000000011000000100101000; // d_in = 4.501953, d_out = 1.504511
				11'd1794: d_out <= 32'b00000000000000011000000101000100; // d_in = 4.503906, d_out = 1.504945
				11'd1795: d_out <= 32'b00000000000000011000000101100000; // d_in = 4.505859, d_out = 1.505379
				11'd1796: d_out <= 32'b00000000000000011000000101111101; // d_in = 4.507812, d_out = 1.505812
				11'd1797: d_out <= 32'b00000000000000011000000110011001; // d_in = 4.509766, d_out = 1.506245
				11'd1798: d_out <= 32'b00000000000000011000000110110110; // d_in = 4.511719, d_out = 1.506678
				11'd1799: d_out <= 32'b00000000000000011000000111010010; // d_in = 4.513672, d_out = 1.507111
				11'd1800: d_out <= 32'b00000000000000011000000111101110; // d_in = 4.515625, d_out = 1.507544
				11'd1801: d_out <= 32'b00000000000000011000001000001011; // d_in = 4.517578, d_out = 1.507976
				11'd1802: d_out <= 32'b00000000000000011000001000100111; // d_in = 4.519531, d_out = 1.508408
				11'd1803: d_out <= 32'b00000000000000011000001001000011; // d_in = 4.521484, d_out = 1.508840
				11'd1804: d_out <= 32'b00000000000000011000001001100000; // d_in = 4.523438, d_out = 1.509272
				11'd1805: d_out <= 32'b00000000000000011000001001111100; // d_in = 4.525391, d_out = 1.509704
				11'd1806: d_out <= 32'b00000000000000011000001010011000; // d_in = 4.527344, d_out = 1.510135
				11'd1807: d_out <= 32'b00000000000000011000001010110101; // d_in = 4.529297, d_out = 1.510567
				11'd1808: d_out <= 32'b00000000000000011000001011010001; // d_in = 4.531250, d_out = 1.510998
				11'd1809: d_out <= 32'b00000000000000011000001011101101; // d_in = 4.533203, d_out = 1.511429
				11'd1810: d_out <= 32'b00000000000000011000001100001001; // d_in = 4.535156, d_out = 1.511860
				11'd1811: d_out <= 32'b00000000000000011000001100100101; // d_in = 4.537109, d_out = 1.512290
				11'd1812: d_out <= 32'b00000000000000011000001101000010; // d_in = 4.539062, d_out = 1.512720
				11'd1813: d_out <= 32'b00000000000000011000001101011110; // d_in = 4.541016, d_out = 1.513151
				11'd1814: d_out <= 32'b00000000000000011000001101111010; // d_in = 4.542969, d_out = 1.513581
				11'd1815: d_out <= 32'b00000000000000011000001110010110; // d_in = 4.544922, d_out = 1.514011
				11'd1816: d_out <= 32'b00000000000000011000001110110010; // d_in = 4.546875, d_out = 1.514440
				11'd1817: d_out <= 32'b00000000000000011000001111001110; // d_in = 4.548828, d_out = 1.514870
				11'd1818: d_out <= 32'b00000000000000011000001111101011; // d_in = 4.550781, d_out = 1.515299
				11'd1819: d_out <= 32'b00000000000000011000010000000111; // d_in = 4.552734, d_out = 1.515728
				11'd1820: d_out <= 32'b00000000000000011000010000100011; // d_in = 4.554688, d_out = 1.516157
				11'd1821: d_out <= 32'b00000000000000011000010000111111; // d_in = 4.556641, d_out = 1.516586
				11'd1822: d_out <= 32'b00000000000000011000010001011011; // d_in = 4.558594, d_out = 1.517014
				11'd1823: d_out <= 32'b00000000000000011000010001110111; // d_in = 4.560547, d_out = 1.517443
				11'd1824: d_out <= 32'b00000000000000011000010010010011; // d_in = 4.562500, d_out = 1.517871
				11'd1825: d_out <= 32'b00000000000000011000010010101111; // d_in = 4.564453, d_out = 1.518299
				11'd1826: d_out <= 32'b00000000000000011000010011001011; // d_in = 4.566406, d_out = 1.518727
				11'd1827: d_out <= 32'b00000000000000011000010011100111; // d_in = 4.568359, d_out = 1.519154
				11'd1828: d_out <= 32'b00000000000000011000010100000011; // d_in = 4.570312, d_out = 1.519582
				11'd1829: d_out <= 32'b00000000000000011000010100011111; // d_in = 4.572266, d_out = 1.520009
				11'd1830: d_out <= 32'b00000000000000011000010100111011; // d_in = 4.574219, d_out = 1.520436
				11'd1831: d_out <= 32'b00000000000000011000010101010111; // d_in = 4.576172, d_out = 1.520863
				11'd1832: d_out <= 32'b00000000000000011000010101110011; // d_in = 4.578125, d_out = 1.521290
				11'd1833: d_out <= 32'b00000000000000011000010110001111; // d_in = 4.580078, d_out = 1.521716
				11'd1834: d_out <= 32'b00000000000000011000010110101011; // d_in = 4.582031, d_out = 1.522142
				11'd1835: d_out <= 32'b00000000000000011000010111000111; // d_in = 4.583984, d_out = 1.522569
				11'd1836: d_out <= 32'b00000000000000011000010111100011; // d_in = 4.585938, d_out = 1.522995
				11'd1837: d_out <= 32'b00000000000000011000010111111111; // d_in = 4.587891, d_out = 1.523420
				11'd1838: d_out <= 32'b00000000000000011000011000011011; // d_in = 4.589844, d_out = 1.523846
				11'd1839: d_out <= 32'b00000000000000011000011000110111; // d_in = 4.591797, d_out = 1.524271
				11'd1840: d_out <= 32'b00000000000000011000011001010011; // d_in = 4.593750, d_out = 1.524697
				11'd1841: d_out <= 32'b00000000000000011000011001101110; // d_in = 4.595703, d_out = 1.525122
				11'd1842: d_out <= 32'b00000000000000011000011010001010; // d_in = 4.597656, d_out = 1.525547
				11'd1843: d_out <= 32'b00000000000000011000011010100110; // d_in = 4.599609, d_out = 1.525971
				11'd1844: d_out <= 32'b00000000000000011000011011000010; // d_in = 4.601562, d_out = 1.526396
				11'd1845: d_out <= 32'b00000000000000011000011011011110; // d_in = 4.603516, d_out = 1.526820
				11'd1846: d_out <= 32'b00000000000000011000011011111001; // d_in = 4.605469, d_out = 1.527244
				11'd1847: d_out <= 32'b00000000000000011000011100010101; // d_in = 4.607422, d_out = 1.527668
				11'd1848: d_out <= 32'b00000000000000011000011100110001; // d_in = 4.609375, d_out = 1.528092
				11'd1849: d_out <= 32'b00000000000000011000011101001101; // d_in = 4.611328, d_out = 1.528516
				11'd1850: d_out <= 32'b00000000000000011000011101101001; // d_in = 4.613281, d_out = 1.528939
				11'd1851: d_out <= 32'b00000000000000011000011110000100; // d_in = 4.615234, d_out = 1.529363
				11'd1852: d_out <= 32'b00000000000000011000011110100000; // d_in = 4.617188, d_out = 1.529786
				11'd1853: d_out <= 32'b00000000000000011000011110111100; // d_in = 4.619141, d_out = 1.530209
				11'd1854: d_out <= 32'b00000000000000011000011111010111; // d_in = 4.621094, d_out = 1.530631
				11'd1855: d_out <= 32'b00000000000000011000011111110011; // d_in = 4.623047, d_out = 1.531054
				11'd1856: d_out <= 32'b00000000000000011000100000001111; // d_in = 4.625000, d_out = 1.531476
				11'd1857: d_out <= 32'b00000000000000011000100000101011; // d_in = 4.626953, d_out = 1.531899
				11'd1858: d_out <= 32'b00000000000000011000100001000110; // d_in = 4.628906, d_out = 1.532321
				11'd1859: d_out <= 32'b00000000000000011000100001100010; // d_in = 4.630859, d_out = 1.532742
				11'd1860: d_out <= 32'b00000000000000011000100001111101; // d_in = 4.632812, d_out = 1.533164
				11'd1861: d_out <= 32'b00000000000000011000100010011001; // d_in = 4.634766, d_out = 1.533586
				11'd1862: d_out <= 32'b00000000000000011000100010110101; // d_in = 4.636719, d_out = 1.534007
				11'd1863: d_out <= 32'b00000000000000011000100011010000; // d_in = 4.638672, d_out = 1.534428
				11'd1864: d_out <= 32'b00000000000000011000100011101100; // d_in = 4.640625, d_out = 1.534849
				11'd1865: d_out <= 32'b00000000000000011000100100000111; // d_in = 4.642578, d_out = 1.535270
				11'd1866: d_out <= 32'b00000000000000011000100100100011; // d_in = 4.644531, d_out = 1.535690
				11'd1867: d_out <= 32'b00000000000000011000100100111111; // d_in = 4.646484, d_out = 1.536111
				11'd1868: d_out <= 32'b00000000000000011000100101011010; // d_in = 4.648438, d_out = 1.536531
				11'd1869: d_out <= 32'b00000000000000011000100101110110; // d_in = 4.650391, d_out = 1.536951
				11'd1870: d_out <= 32'b00000000000000011000100110010001; // d_in = 4.652344, d_out = 1.537371
				11'd1871: d_out <= 32'b00000000000000011000100110101101; // d_in = 4.654297, d_out = 1.537791
				11'd1872: d_out <= 32'b00000000000000011000100111001000; // d_in = 4.656250, d_out = 1.538210
				11'd1873: d_out <= 32'b00000000000000011000100111100100; // d_in = 4.658203, d_out = 1.538630
				11'd1874: d_out <= 32'b00000000000000011000100111111111; // d_in = 4.660156, d_out = 1.539049
				11'd1875: d_out <= 32'b00000000000000011000101000011011; // d_in = 4.662109, d_out = 1.539468
				11'd1876: d_out <= 32'b00000000000000011000101000110110; // d_in = 4.664062, d_out = 1.539887
				11'd1877: d_out <= 32'b00000000000000011000101001010001; // d_in = 4.666016, d_out = 1.540306
				11'd1878: d_out <= 32'b00000000000000011000101001101101; // d_in = 4.667969, d_out = 1.540724
				11'd1879: d_out <= 32'b00000000000000011000101010001000; // d_in = 4.669922, d_out = 1.541142
				11'd1880: d_out <= 32'b00000000000000011000101010100100; // d_in = 4.671875, d_out = 1.541560
				11'd1881: d_out <= 32'b00000000000000011000101010111111; // d_in = 4.673828, d_out = 1.541978
				11'd1882: d_out <= 32'b00000000000000011000101011011010; // d_in = 4.675781, d_out = 1.542396
				11'd1883: d_out <= 32'b00000000000000011000101011110110; // d_in = 4.677734, d_out = 1.542814
				11'd1884: d_out <= 32'b00000000000000011000101100010001; // d_in = 4.679688, d_out = 1.543231
				11'd1885: d_out <= 32'b00000000000000011000101100101101; // d_in = 4.681641, d_out = 1.543649
				11'd1886: d_out <= 32'b00000000000000011000101101001000; // d_in = 4.683594, d_out = 1.544066
				11'd1887: d_out <= 32'b00000000000000011000101101100011; // d_in = 4.685547, d_out = 1.544483
				11'd1888: d_out <= 32'b00000000000000011000101101111111; // d_in = 4.687500, d_out = 1.544899
				11'd1889: d_out <= 32'b00000000000000011000101110011010; // d_in = 4.689453, d_out = 1.545316
				11'd1890: d_out <= 32'b00000000000000011000101110110101; // d_in = 4.691406, d_out = 1.545732
				11'd1891: d_out <= 32'b00000000000000011000101111010000; // d_in = 4.693359, d_out = 1.546149
				11'd1892: d_out <= 32'b00000000000000011000101111101100; // d_in = 4.695312, d_out = 1.546565
				11'd1893: d_out <= 32'b00000000000000011000110000000111; // d_in = 4.697266, d_out = 1.546981
				11'd1894: d_out <= 32'b00000000000000011000110000100010; // d_in = 4.699219, d_out = 1.547396
				11'd1895: d_out <= 32'b00000000000000011000110000111101; // d_in = 4.701172, d_out = 1.547812
				11'd1896: d_out <= 32'b00000000000000011000110001011001; // d_in = 4.703125, d_out = 1.548227
				11'd1897: d_out <= 32'b00000000000000011000110001110100; // d_in = 4.705078, d_out = 1.548642
				11'd1898: d_out <= 32'b00000000000000011000110010001111; // d_in = 4.707031, d_out = 1.549057
				11'd1899: d_out <= 32'b00000000000000011000110010101010; // d_in = 4.708984, d_out = 1.549472
				11'd1900: d_out <= 32'b00000000000000011000110011000101; // d_in = 4.710938, d_out = 1.549887
				11'd1901: d_out <= 32'b00000000000000011000110011100001; // d_in = 4.712891, d_out = 1.550301
				11'd1902: d_out <= 32'b00000000000000011000110011111100; // d_in = 4.714844, d_out = 1.550716
				11'd1903: d_out <= 32'b00000000000000011000110100010111; // d_in = 4.716797, d_out = 1.551130
				11'd1904: d_out <= 32'b00000000000000011000110100110010; // d_in = 4.718750, d_out = 1.551544
				11'd1905: d_out <= 32'b00000000000000011000110101001101; // d_in = 4.720703, d_out = 1.551958
				11'd1906: d_out <= 32'b00000000000000011000110101101000; // d_in = 4.722656, d_out = 1.552371
				11'd1907: d_out <= 32'b00000000000000011000110110000011; // d_in = 4.724609, d_out = 1.552785
				11'd1908: d_out <= 32'b00000000000000011000110110011110; // d_in = 4.726562, d_out = 1.553198
				11'd1909: d_out <= 32'b00000000000000011000110110111001; // d_in = 4.728516, d_out = 1.553611
				11'd1910: d_out <= 32'b00000000000000011000110111010101; // d_in = 4.730469, d_out = 1.554024
				11'd1911: d_out <= 32'b00000000000000011000110111110000; // d_in = 4.732422, d_out = 1.554437
				11'd1912: d_out <= 32'b00000000000000011000111000001011; // d_in = 4.734375, d_out = 1.554850
				11'd1913: d_out <= 32'b00000000000000011000111000100110; // d_in = 4.736328, d_out = 1.555262
				11'd1914: d_out <= 32'b00000000000000011000111001000001; // d_in = 4.738281, d_out = 1.555674
				11'd1915: d_out <= 32'b00000000000000011000111001011100; // d_in = 4.740234, d_out = 1.556087
				11'd1916: d_out <= 32'b00000000000000011000111001110111; // d_in = 4.742188, d_out = 1.556499
				11'd1917: d_out <= 32'b00000000000000011000111010010010; // d_in = 4.744141, d_out = 1.556910
				11'd1918: d_out <= 32'b00000000000000011000111010101101; // d_in = 4.746094, d_out = 1.557322
				11'd1919: d_out <= 32'b00000000000000011000111011001000; // d_in = 4.748047, d_out = 1.557733
				11'd1920: d_out <= 32'b00000000000000011000111011100011; // d_in = 4.750000, d_out = 1.558145
				11'd1921: d_out <= 32'b00000000000000011000111011111110; // d_in = 4.751953, d_out = 1.558556
				11'd1922: d_out <= 32'b00000000000000011000111100011000; // d_in = 4.753906, d_out = 1.558967
				11'd1923: d_out <= 32'b00000000000000011000111100110011; // d_in = 4.755859, d_out = 1.559377
				11'd1924: d_out <= 32'b00000000000000011000111101001110; // d_in = 4.757812, d_out = 1.559788
				11'd1925: d_out <= 32'b00000000000000011000111101101001; // d_in = 4.759766, d_out = 1.560198
				11'd1926: d_out <= 32'b00000000000000011000111110000100; // d_in = 4.761719, d_out = 1.560609
				11'd1927: d_out <= 32'b00000000000000011000111110011111; // d_in = 4.763672, d_out = 1.561019
				11'd1928: d_out <= 32'b00000000000000011000111110111010; // d_in = 4.765625, d_out = 1.561429
				11'd1929: d_out <= 32'b00000000000000011000111111010101; // d_in = 4.767578, d_out = 1.561838
				11'd1930: d_out <= 32'b00000000000000011000111111101111; // d_in = 4.769531, d_out = 1.562248
				11'd1931: d_out <= 32'b00000000000000011001000000001010; // d_in = 4.771484, d_out = 1.562657
				11'd1932: d_out <= 32'b00000000000000011001000000100101; // d_in = 4.773438, d_out = 1.563067
				11'd1933: d_out <= 32'b00000000000000011001000001000000; // d_in = 4.775391, d_out = 1.563476
				11'd1934: d_out <= 32'b00000000000000011001000001011011; // d_in = 4.777344, d_out = 1.563885
				11'd1935: d_out <= 32'b00000000000000011001000001110110; // d_in = 4.779297, d_out = 1.564293
				11'd1936: d_out <= 32'b00000000000000011001000010010000; // d_in = 4.781250, d_out = 1.564702
				11'd1937: d_out <= 32'b00000000000000011001000010101011; // d_in = 4.783203, d_out = 1.565110
				11'd1938: d_out <= 32'b00000000000000011001000011000110; // d_in = 4.785156, d_out = 1.565519
				11'd1939: d_out <= 32'b00000000000000011001000011100001; // d_in = 4.787109, d_out = 1.565927
				11'd1940: d_out <= 32'b00000000000000011001000011111011; // d_in = 4.789062, d_out = 1.566335
				11'd1941: d_out <= 32'b00000000000000011001000100010110; // d_in = 4.791016, d_out = 1.566742
				11'd1942: d_out <= 32'b00000000000000011001000100110001; // d_in = 4.792969, d_out = 1.567150
				11'd1943: d_out <= 32'b00000000000000011001000101001011; // d_in = 4.794922, d_out = 1.567557
				11'd1944: d_out <= 32'b00000000000000011001000101100110; // d_in = 4.796875, d_out = 1.567965
				11'd1945: d_out <= 32'b00000000000000011001000110000001; // d_in = 4.798828, d_out = 1.568372
				11'd1946: d_out <= 32'b00000000000000011001000110011011; // d_in = 4.800781, d_out = 1.568779
				11'd1947: d_out <= 32'b00000000000000011001000110110110; // d_in = 4.802734, d_out = 1.569185
				11'd1948: d_out <= 32'b00000000000000011001000111010001; // d_in = 4.804688, d_out = 1.569592
				11'd1949: d_out <= 32'b00000000000000011001000111101011; // d_in = 4.806641, d_out = 1.569998
				11'd1950: d_out <= 32'b00000000000000011001001000000110; // d_in = 4.808594, d_out = 1.570405
				11'd1951: d_out <= 32'b00000000000000011001001000100001; // d_in = 4.810547, d_out = 1.570811
				11'd1952: d_out <= 32'b00000000000000011001001000111011; // d_in = 4.812500, d_out = 1.571217
				11'd1953: d_out <= 32'b00000000000000011001001001010110; // d_in = 4.814453, d_out = 1.571622
				11'd1954: d_out <= 32'b00000000000000011001001001110000; // d_in = 4.816406, d_out = 1.572028
				11'd1955: d_out <= 32'b00000000000000011001001010001011; // d_in = 4.818359, d_out = 1.572433
				11'd1956: d_out <= 32'b00000000000000011001001010100110; // d_in = 4.820312, d_out = 1.572839
				11'd1957: d_out <= 32'b00000000000000011001001011000000; // d_in = 4.822266, d_out = 1.573244
				11'd1958: d_out <= 32'b00000000000000011001001011011011; // d_in = 4.824219, d_out = 1.573649
				11'd1959: d_out <= 32'b00000000000000011001001011110101; // d_in = 4.826172, d_out = 1.574054
				11'd1960: d_out <= 32'b00000000000000011001001100010000; // d_in = 4.828125, d_out = 1.574458
				11'd1961: d_out <= 32'b00000000000000011001001100101010; // d_in = 4.830078, d_out = 1.574863
				11'd1962: d_out <= 32'b00000000000000011001001101000101; // d_in = 4.832031, d_out = 1.575267
				11'd1963: d_out <= 32'b00000000000000011001001101011111; // d_in = 4.833984, d_out = 1.575671
				11'd1964: d_out <= 32'b00000000000000011001001101111010; // d_in = 4.835938, d_out = 1.576075
				11'd1965: d_out <= 32'b00000000000000011001001110010100; // d_in = 4.837891, d_out = 1.576479
				11'd1966: d_out <= 32'b00000000000000011001001110101111; // d_in = 4.839844, d_out = 1.576882
				11'd1967: d_out <= 32'b00000000000000011001001111001001; // d_in = 4.841797, d_out = 1.577286
				11'd1968: d_out <= 32'b00000000000000011001001111100011; // d_in = 4.843750, d_out = 1.577689
				11'd1969: d_out <= 32'b00000000000000011001001111111110; // d_in = 4.845703, d_out = 1.578092
				11'd1970: d_out <= 32'b00000000000000011001010000011000; // d_in = 4.847656, d_out = 1.578495
				11'd1971: d_out <= 32'b00000000000000011001010000110011; // d_in = 4.849609, d_out = 1.578898
				11'd1972: d_out <= 32'b00000000000000011001010001001101; // d_in = 4.851562, d_out = 1.579301
				11'd1973: d_out <= 32'b00000000000000011001010001100111; // d_in = 4.853516, d_out = 1.579703
				11'd1974: d_out <= 32'b00000000000000011001010010000010; // d_in = 4.855469, d_out = 1.580106
				11'd1975: d_out <= 32'b00000000000000011001010010011100; // d_in = 4.857422, d_out = 1.580508
				11'd1976: d_out <= 32'b00000000000000011001010010110111; // d_in = 4.859375, d_out = 1.580910
				11'd1977: d_out <= 32'b00000000000000011001010011010001; // d_in = 4.861328, d_out = 1.581312
				11'd1978: d_out <= 32'b00000000000000011001010011101011; // d_in = 4.863281, d_out = 1.581713
				11'd1979: d_out <= 32'b00000000000000011001010100000101; // d_in = 4.865234, d_out = 1.582115
				11'd1980: d_out <= 32'b00000000000000011001010100100000; // d_in = 4.867188, d_out = 1.582516
				11'd1981: d_out <= 32'b00000000000000011001010100111010; // d_in = 4.869141, d_out = 1.582917
				11'd1982: d_out <= 32'b00000000000000011001010101010100; // d_in = 4.871094, d_out = 1.583319
				11'd1983: d_out <= 32'b00000000000000011001010101101111; // d_in = 4.873047, d_out = 1.583719
				11'd1984: d_out <= 32'b00000000000000011001010110001001; // d_in = 4.875000, d_out = 1.584120
				11'd1985: d_out <= 32'b00000000000000011001010110100011; // d_in = 4.876953, d_out = 1.584521
				11'd1986: d_out <= 32'b00000000000000011001010110111101; // d_in = 4.878906, d_out = 1.584921
				11'd1987: d_out <= 32'b00000000000000011001010111011000; // d_in = 4.880859, d_out = 1.585321
				11'd1988: d_out <= 32'b00000000000000011001010111110010; // d_in = 4.882812, d_out = 1.585721
				11'd1989: d_out <= 32'b00000000000000011001011000001100; // d_in = 4.884766, d_out = 1.586121
				11'd1990: d_out <= 32'b00000000000000011001011000100110; // d_in = 4.886719, d_out = 1.586521
				11'd1991: d_out <= 32'b00000000000000011001011001000000; // d_in = 4.888672, d_out = 1.586921
				11'd1992: d_out <= 32'b00000000000000011001011001011011; // d_in = 4.890625, d_out = 1.587320
				11'd1993: d_out <= 32'b00000000000000011001011001110101; // d_in = 4.892578, d_out = 1.587719
				11'd1994: d_out <= 32'b00000000000000011001011010001111; // d_in = 4.894531, d_out = 1.588119
				11'd1995: d_out <= 32'b00000000000000011001011010101001; // d_in = 4.896484, d_out = 1.588517
				11'd1996: d_out <= 32'b00000000000000011001011011000011; // d_in = 4.898438, d_out = 1.588916
				11'd1997: d_out <= 32'b00000000000000011001011011011101; // d_in = 4.900391, d_out = 1.589315
				11'd1998: d_out <= 32'b00000000000000011001011011110111; // d_in = 4.902344, d_out = 1.589713
				11'd1999: d_out <= 32'b00000000000000011001011100010010; // d_in = 4.904297, d_out = 1.590112
				11'd2000: d_out <= 32'b00000000000000011001011100101100; // d_in = 4.906250, d_out = 1.590510
				11'd2001: d_out <= 32'b00000000000000011001011101000110; // d_in = 4.908203, d_out = 1.590908
				11'd2002: d_out <= 32'b00000000000000011001011101100000; // d_in = 4.910156, d_out = 1.591306
				11'd2003: d_out <= 32'b00000000000000011001011101111010; // d_in = 4.912109, d_out = 1.591703
				11'd2004: d_out <= 32'b00000000000000011001011110010100; // d_in = 4.914062, d_out = 1.592101
				11'd2005: d_out <= 32'b00000000000000011001011110101110; // d_in = 4.916016, d_out = 1.592498
				11'd2006: d_out <= 32'b00000000000000011001011111001000; // d_in = 4.917969, d_out = 1.592896
				11'd2007: d_out <= 32'b00000000000000011001011111100010; // d_in = 4.919922, d_out = 1.593293
				11'd2008: d_out <= 32'b00000000000000011001011111111100; // d_in = 4.921875, d_out = 1.593690
				11'd2009: d_out <= 32'b00000000000000011001100000010110; // d_in = 4.923828, d_out = 1.594086
				11'd2010: d_out <= 32'b00000000000000011001100000110000; // d_in = 4.925781, d_out = 1.594483
				11'd2011: d_out <= 32'b00000000000000011001100001001010; // d_in = 4.927734, d_out = 1.594879
				11'd2012: d_out <= 32'b00000000000000011001100001100100; // d_in = 4.929688, d_out = 1.595276
				11'd2013: d_out <= 32'b00000000000000011001100001111110; // d_in = 4.931641, d_out = 1.595672
				11'd2014: d_out <= 32'b00000000000000011001100010011000; // d_in = 4.933594, d_out = 1.596068
				11'd2015: d_out <= 32'b00000000000000011001100010110010; // d_in = 4.935547, d_out = 1.596463
				11'd2016: d_out <= 32'b00000000000000011001100011001100; // d_in = 4.937500, d_out = 1.596859
				11'd2017: d_out <= 32'b00000000000000011001100011100110; // d_in = 4.939453, d_out = 1.597255
				11'd2018: d_out <= 32'b00000000000000011001100100000000; // d_in = 4.941406, d_out = 1.597650
				11'd2019: d_out <= 32'b00000000000000011001100100011001; // d_in = 4.943359, d_out = 1.598045
				11'd2020: d_out <= 32'b00000000000000011001100100110011; // d_in = 4.945312, d_out = 1.598440
				11'd2021: d_out <= 32'b00000000000000011001100101001101; // d_in = 4.947266, d_out = 1.598835
				11'd2022: d_out <= 32'b00000000000000011001100101100111; // d_in = 4.949219, d_out = 1.599230
				11'd2023: d_out <= 32'b00000000000000011001100110000001; // d_in = 4.951172, d_out = 1.599624
				11'd2024: d_out <= 32'b00000000000000011001100110011011; // d_in = 4.953125, d_out = 1.600019
				11'd2025: d_out <= 32'b00000000000000011001100110110101; // d_in = 4.955078, d_out = 1.600413
				11'd2026: d_out <= 32'b00000000000000011001100111001110; // d_in = 4.957031, d_out = 1.600807
				11'd2027: d_out <= 32'b00000000000000011001100111101000; // d_in = 4.958984, d_out = 1.601201
				11'd2028: d_out <= 32'b00000000000000011001101000000010; // d_in = 4.960938, d_out = 1.601595
				11'd2029: d_out <= 32'b00000000000000011001101000011100; // d_in = 4.962891, d_out = 1.601988
				11'd2030: d_out <= 32'b00000000000000011001101000110110; // d_in = 4.964844, d_out = 1.602382
				11'd2031: d_out <= 32'b00000000000000011001101001001111; // d_in = 4.966797, d_out = 1.602775
				11'd2032: d_out <= 32'b00000000000000011001101001101001; // d_in = 4.968750, d_out = 1.603168
				11'd2033: d_out <= 32'b00000000000000011001101010000011; // d_in = 4.970703, d_out = 1.603561
				11'd2034: d_out <= 32'b00000000000000011001101010011101; // d_in = 4.972656, d_out = 1.603954
				11'd2035: d_out <= 32'b00000000000000011001101010110110; // d_in = 4.974609, d_out = 1.604347
				11'd2036: d_out <= 32'b00000000000000011001101011010000; // d_in = 4.976562, d_out = 1.604739
				11'd2037: d_out <= 32'b00000000000000011001101011101010; // d_in = 4.978516, d_out = 1.605132
				11'd2038: d_out <= 32'b00000000000000011001101100000100; // d_in = 4.980469, d_out = 1.605524
				11'd2039: d_out <= 32'b00000000000000011001101100011101; // d_in = 4.982422, d_out = 1.605916
				11'd2040: d_out <= 32'b00000000000000011001101100110111; // d_in = 4.984375, d_out = 1.606308
				11'd2041: d_out <= 32'b00000000000000011001101101010001; // d_in = 4.986328, d_out = 1.606700
				11'd2042: d_out <= 32'b00000000000000011001101101101010; // d_in = 4.988281, d_out = 1.607091
				11'd2043: d_out <= 32'b00000000000000011001101110000100; // d_in = 4.990234, d_out = 1.607483
				11'd2044: d_out <= 32'b00000000000000011001101110011110; // d_in = 4.992188, d_out = 1.607874
				11'd2045: d_out <= 32'b00000000000000011001101110110111; // d_in = 4.994141, d_out = 1.608265
				11'd2046: d_out <= 32'b00000000000000011001101111010001; // d_in = 4.996094, d_out = 1.608656
				11'd2047: d_out <= 32'b00000000000000011001101111101011; // d_in = 4.998047, d_out = 1.609047
			endcase
		end
	address_gen u_address_gen(d_in, addr);
endmodule
module address_gen(d_in, addr);
	input  [31:0] d_in;
	output [10:0] addr;

	wire   [1:0] diff;
	assign diff = d_in[18:16] - 3'd1;
	assign addr = {diff, d_in[15:7]};
endmodule
