/*----------------------------------------------------------------------------
  Copyright (c) 2004 Aoki laboratory. All rights reserved.

  Top module: multiplier_32b

  Number system: 2's complement
  Multiplicand length: 32
  Multiplier length: 32
  Partial product generation: Simple PPG
  Partial product accumulation: Wallace tree
  Final stage addition: Kogge-Stone adder
----------------------------------------------------------------------------*/
// Modified by: Amir Yazdanbakhsh
// Email: a.yazdanbakhsh@gatech.edu

`timescale 1ns/1ps

module TCDECON_31_0(TOP, R, I);
  output [30:0] R;
  output [31:31] TOP;
  input [31:0] I;
  assign TOP[31] = I[31];
  assign R[0] = I[0];
  assign R[1] = I[1];
  assign R[2] = I[2];
  assign R[3] = I[3];
  assign R[4] = I[4];
  assign R[5] = I[5];
  assign R[6] = I[6];
  assign R[7] = I[7];
  assign R[8] = I[8];
  assign R[9] = I[9];
  assign R[10] = I[10];
  assign R[11] = I[11];
  assign R[12] = I[12];
  assign R[13] = I[13];
  assign R[14] = I[14];
  assign R[15] = I[15];
  assign R[16] = I[16];
  assign R[17] = I[17];
  assign R[18] = I[18];
  assign R[19] = I[19];
  assign R[20] = I[20];
  assign R[21] = I[21];
  assign R[22] = I[22];
  assign R[23] = I[23];
  assign R[24] = I[24];
  assign R[25] = I[25];
  assign R[26] = I[26];
  assign R[27] = I[27];
  assign R[28] = I[28];
  assign R[29] = I[29];
  assign R[30] = I[30];
endmodule

module UB1BPPG_0_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_0(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_31(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_1(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_32(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_2(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_33(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_3(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_34(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_4(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_35(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_5(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_36(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_6(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_37(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_7(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_38(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_8(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_39(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_9(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_40(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_10(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_41(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_11(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_42(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_12(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_43(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_13(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_44(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_14(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_45(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_15(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_46(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_16(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_47(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_17(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_48(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_18(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_49(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_19(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_50(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_20(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_51(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_21(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_52(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_22(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_53(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_23(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_54(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_24(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_55(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_25(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_56(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_26(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_57(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_27(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_58(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_28(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_59(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_29(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_60(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UB1BPPG_0_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_1_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_2_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_3_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_4_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_5_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_6_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_7_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_8_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_9_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_10_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_11_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_12_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_13_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_14_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_15_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_16_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_17_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_18_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_19_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_20_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_21_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_22_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_23_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_24_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_25_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_26_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_27_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_28_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_29_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UB1BPPG_30_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NU1BPPG_31_30(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUBUB1CON_61(O, I);
  output O;
  input I;
  assign O = ~ I;
endmodule

module UN1BPPG_0_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_1_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_2_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_3_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_4_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_5_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_6_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_7_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_8_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_9_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_10_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_11_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_12_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_13_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_14_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_15_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_16_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_17_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_18_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_19_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_20_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_21_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_22_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_23_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_24_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_25_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_26_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_27_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_28_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_29_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UN1BPPG_30_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module NUB1BPPG_31_31(O, IN1, IN2);
  output O;
  input IN1;
  input IN2;
  assign O = IN1 & IN2;
endmodule

module UBOne_32(O);
  output O;
  assign O = 1;
endmodule

module UB1DCON_32(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_1(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_2(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_3(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_4(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_5(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_6(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_7(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_8(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_9(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_10(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_11(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_12(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_13(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_14(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_15(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_16(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_17(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_18(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_19(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_20(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_21(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_22(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_23(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_24(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_25(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_26(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_27(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_28(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_29(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_30(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_31(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_32(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_33(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_4(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_33(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_34(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_35(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_36(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_7(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_35(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_36(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_37(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_38(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_39(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_10(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_38(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_39(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_40(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_41(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_42(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_2(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_34(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_35(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_6(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_37(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_39(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_11(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_41(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_42(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UB1DCON_43(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_14(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_43(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_44(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_45(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_46(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_17(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_45(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_46(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_47(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_48(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_49(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_20(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_48(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_49(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_50(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_51(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_52(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_23(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_51(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_52(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_53(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_54(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_55(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_26(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_54(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_55(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_56(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_57(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_58(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_29(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_57(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_58(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_59(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_60(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_61(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_3(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_36(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_37(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_38(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_9(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_42(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_43(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_15(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_47(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_48(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_19(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_50(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_52(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_24(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_56(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_57(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_28(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_59(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_61(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_5(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_40(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_41(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_13(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_46(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_47(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_21(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_53(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_54(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_27(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_58(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_62(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_8(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_44(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_45(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_18(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_49(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_30(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBFA_60(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_61(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBFA_62(C, S, X, Y, Z);
  output C;
  output S;
  input X;
  input Y;
  input Z;
  assign C = ( X & Y ) | ( Y & Z ) | ( Z & X );
  assign S = X ^ Y ^ Z;
endmodule

module UBHA_12(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_50(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_51(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_53(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_25(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_56(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_62(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_63(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_16(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_55(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UB1DCON_59(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UB1DCON_60(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBHA_22(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBHA_63(C, S, X, Y);
  output C;
  output S;
  input X;
  input Y;
  assign C = X & Y;
  assign S = X ^ Y;
endmodule

module UBZero_64_64(O);
  output [64:64] O;
  assign O[64] = 0;
endmodule

module GPGenerator(Go, Po, A, B);
  output Go;
  output Po;
  input A;
  input B;
  assign Go = A & B;
  assign Po = A ^ B;
endmodule

module CarryOperator(Go, Po, Gi1, Pi1, Gi2, Pi2);
  output Go;
  output Po;
  input Gi1;
  input Gi2;
  input Pi1;
  input Pi2;
  assign Go = Gi1 | ( Gi2 & Pi1 );
  assign Po = Pi1 & Pi2;
endmodule

module UBPriKSA_64_9(S, X, Y, Cin);
  output [65:9] S;
  input Cin;
  input [64:9] X;
  input [64:9] Y;
  wire [64:9] G0;
  wire [64:9] G1;
  wire [64:9] G2;
  wire [64:9] G3;
  wire [64:9] G4;
  wire [64:9] G5;
  wire [64:9] G6;
  wire [64:9] P0;
  wire [64:9] P1;
  wire [64:9] P2;
  wire [64:9] P3;
  wire [64:9] P4;
  wire [64:9] P5;
  wire [64:9] P6;
  assign P1[9] = P0[9];
  assign G1[9] = G0[9];
  assign P2[9] = P1[9];
  assign G2[9] = G1[9];
  assign P2[10] = P1[10];
  assign G2[10] = G1[10];
  assign P3[9] = P2[9];
  assign G3[9] = G2[9];
  assign P3[10] = P2[10];
  assign G3[10] = G2[10];
  assign P3[11] = P2[11];
  assign G3[11] = G2[11];
  assign P3[12] = P2[12];
  assign G3[12] = G2[12];
  assign P4[9] = P3[9];
  assign G4[9] = G3[9];
  assign P4[10] = P3[10];
  assign G4[10] = G3[10];
  assign P4[11] = P3[11];
  assign G4[11] = G3[11];
  assign P4[12] = P3[12];
  assign G4[12] = G3[12];
  assign P4[13] = P3[13];
  assign G4[13] = G3[13];
  assign P4[14] = P3[14];
  assign G4[14] = G3[14];
  assign P4[15] = P3[15];
  assign G4[15] = G3[15];
  assign P4[16] = P3[16];
  assign G4[16] = G3[16];
  assign P5[9] = P4[9];
  assign G5[9] = G4[9];
  assign P5[10] = P4[10];
  assign G5[10] = G4[10];
  assign P5[11] = P4[11];
  assign G5[11] = G4[11];
  assign P5[12] = P4[12];
  assign G5[12] = G4[12];
  assign P5[13] = P4[13];
  assign G5[13] = G4[13];
  assign P5[14] = P4[14];
  assign G5[14] = G4[14];
  assign P5[15] = P4[15];
  assign G5[15] = G4[15];
  assign P5[16] = P4[16];
  assign G5[16] = G4[16];
  assign P5[17] = P4[17];
  assign G5[17] = G4[17];
  assign P5[18] = P4[18];
  assign G5[18] = G4[18];
  assign P5[19] = P4[19];
  assign G5[19] = G4[19];
  assign P5[20] = P4[20];
  assign G5[20] = G4[20];
  assign P5[21] = P4[21];
  assign G5[21] = G4[21];
  assign P5[22] = P4[22];
  assign G5[22] = G4[22];
  assign P5[23] = P4[23];
  assign G5[23] = G4[23];
  assign P5[24] = P4[24];
  assign G5[24] = G4[24];
  assign P6[9] = P5[9];
  assign G6[9] = G5[9];
  assign P6[10] = P5[10];
  assign G6[10] = G5[10];
  assign P6[11] = P5[11];
  assign G6[11] = G5[11];
  assign P6[12] = P5[12];
  assign G6[12] = G5[12];
  assign P6[13] = P5[13];
  assign G6[13] = G5[13];
  assign P6[14] = P5[14];
  assign G6[14] = G5[14];
  assign P6[15] = P5[15];
  assign G6[15] = G5[15];
  assign P6[16] = P5[16];
  assign G6[16] = G5[16];
  assign P6[17] = P5[17];
  assign G6[17] = G5[17];
  assign P6[18] = P5[18];
  assign G6[18] = G5[18];
  assign P6[19] = P5[19];
  assign G6[19] = G5[19];
  assign P6[20] = P5[20];
  assign G6[20] = G5[20];
  assign P6[21] = P5[21];
  assign G6[21] = G5[21];
  assign P6[22] = P5[22];
  assign G6[22] = G5[22];
  assign P6[23] = P5[23];
  assign G6[23] = G5[23];
  assign P6[24] = P5[24];
  assign G6[24] = G5[24];
  assign P6[25] = P5[25];
  assign G6[25] = G5[25];
  assign P6[26] = P5[26];
  assign G6[26] = G5[26];
  assign P6[27] = P5[27];
  assign G6[27] = G5[27];
  assign P6[28] = P5[28];
  assign G6[28] = G5[28];
  assign P6[29] = P5[29];
  assign G6[29] = G5[29];
  assign P6[30] = P5[30];
  assign G6[30] = G5[30];
  assign P6[31] = P5[31];
  assign G6[31] = G5[31];
  assign P6[32] = P5[32];
  assign G6[32] = G5[32];
  assign P6[33] = P5[33];
  assign G6[33] = G5[33];
  assign P6[34] = P5[34];
  assign G6[34] = G5[34];
  assign P6[35] = P5[35];
  assign G6[35] = G5[35];
  assign P6[36] = P5[36];
  assign G6[36] = G5[36];
  assign P6[37] = P5[37];
  assign G6[37] = G5[37];
  assign P6[38] = P5[38];
  assign G6[38] = G5[38];
  assign P6[39] = P5[39];
  assign G6[39] = G5[39];
  assign P6[40] = P5[40];
  assign G6[40] = G5[40];
  assign S[9] = Cin ^ P0[9];
  assign S[10] = ( G6[9] | ( P6[9] & Cin ) ) ^ P0[10];
  assign S[11] = ( G6[10] | ( P6[10] & Cin ) ) ^ P0[11];
  assign S[12] = ( G6[11] | ( P6[11] & Cin ) ) ^ P0[12];
  assign S[13] = ( G6[12] | ( P6[12] & Cin ) ) ^ P0[13];
  assign S[14] = ( G6[13] | ( P6[13] & Cin ) ) ^ P0[14];
  assign S[15] = ( G6[14] | ( P6[14] & Cin ) ) ^ P0[15];
  assign S[16] = ( G6[15] | ( P6[15] & Cin ) ) ^ P0[16];
  assign S[17] = ( G6[16] | ( P6[16] & Cin ) ) ^ P0[17];
  assign S[18] = ( G6[17] | ( P6[17] & Cin ) ) ^ P0[18];
  assign S[19] = ( G6[18] | ( P6[18] & Cin ) ) ^ P0[19];
  assign S[20] = ( G6[19] | ( P6[19] & Cin ) ) ^ P0[20];
  assign S[21] = ( G6[20] | ( P6[20] & Cin ) ) ^ P0[21];
  assign S[22] = ( G6[21] | ( P6[21] & Cin ) ) ^ P0[22];
  assign S[23] = ( G6[22] | ( P6[22] & Cin ) ) ^ P0[23];
  assign S[24] = ( G6[23] | ( P6[23] & Cin ) ) ^ P0[24];
  assign S[25] = ( G6[24] | ( P6[24] & Cin ) ) ^ P0[25];
  assign S[26] = ( G6[25] | ( P6[25] & Cin ) ) ^ P0[26];
  assign S[27] = ( G6[26] | ( P6[26] & Cin ) ) ^ P0[27];
  assign S[28] = ( G6[27] | ( P6[27] & Cin ) ) ^ P0[28];
  assign S[29] = ( G6[28] | ( P6[28] & Cin ) ) ^ P0[29];
  assign S[30] = ( G6[29] | ( P6[29] & Cin ) ) ^ P0[30];
  assign S[31] = ( G6[30] | ( P6[30] & Cin ) ) ^ P0[31];
  assign S[32] = ( G6[31] | ( P6[31] & Cin ) ) ^ P0[32];
  assign S[33] = ( G6[32] | ( P6[32] & Cin ) ) ^ P0[33];
  assign S[34] = ( G6[33] | ( P6[33] & Cin ) ) ^ P0[34];
  assign S[35] = ( G6[34] | ( P6[34] & Cin ) ) ^ P0[35];
  assign S[36] = ( G6[35] | ( P6[35] & Cin ) ) ^ P0[36];
  assign S[37] = ( G6[36] | ( P6[36] & Cin ) ) ^ P0[37];
  assign S[38] = ( G6[37] | ( P6[37] & Cin ) ) ^ P0[38];
  assign S[39] = ( G6[38] | ( P6[38] & Cin ) ) ^ P0[39];
  assign S[40] = ( G6[39] | ( P6[39] & Cin ) ) ^ P0[40];
  assign S[41] = ( G6[40] | ( P6[40] & Cin ) ) ^ P0[41];
  assign S[42] = ( G6[41] | ( P6[41] & Cin ) ) ^ P0[42];
  assign S[43] = ( G6[42] | ( P6[42] & Cin ) ) ^ P0[43];
  assign S[44] = ( G6[43] | ( P6[43] & Cin ) ) ^ P0[44];
  assign S[45] = ( G6[44] | ( P6[44] & Cin ) ) ^ P0[45];
  assign S[46] = ( G6[45] | ( P6[45] & Cin ) ) ^ P0[46];
  assign S[47] = ( G6[46] | ( P6[46] & Cin ) ) ^ P0[47];
  assign S[48] = ( G6[47] | ( P6[47] & Cin ) ) ^ P0[48];
  assign S[49] = ( G6[48] | ( P6[48] & Cin ) ) ^ P0[49];
  assign S[50] = ( G6[49] | ( P6[49] & Cin ) ) ^ P0[50];
  assign S[51] = ( G6[50] | ( P6[50] & Cin ) ) ^ P0[51];
  assign S[52] = ( G6[51] | ( P6[51] & Cin ) ) ^ P0[52];
  assign S[53] = ( G6[52] | ( P6[52] & Cin ) ) ^ P0[53];
  assign S[54] = ( G6[53] | ( P6[53] & Cin ) ) ^ P0[54];
  assign S[55] = ( G6[54] | ( P6[54] & Cin ) ) ^ P0[55];
  assign S[56] = ( G6[55] | ( P6[55] & Cin ) ) ^ P0[56];
  assign S[57] = ( G6[56] | ( P6[56] & Cin ) ) ^ P0[57];
  assign S[58] = ( G6[57] | ( P6[57] & Cin ) ) ^ P0[58];
  assign S[59] = ( G6[58] | ( P6[58] & Cin ) ) ^ P0[59];
  assign S[60] = ( G6[59] | ( P6[59] & Cin ) ) ^ P0[60];
  assign S[61] = ( G6[60] | ( P6[60] & Cin ) ) ^ P0[61];
  assign S[62] = ( G6[61] | ( P6[61] & Cin ) ) ^ P0[62];
  assign S[63] = ( G6[62] | ( P6[62] & Cin ) ) ^ P0[63];
  assign S[64] = ( G6[63] | ( P6[63] & Cin ) ) ^ P0[64];
  assign S[65] = G6[64] | ( P6[64] & Cin );
  GPGenerator U0 (G0[9], P0[9], X[9], Y[9]);
  GPGenerator U1 (G0[10], P0[10], X[10], Y[10]);
  GPGenerator U2 (G0[11], P0[11], X[11], Y[11]);
  GPGenerator U3 (G0[12], P0[12], X[12], Y[12]);
  GPGenerator U4 (G0[13], P0[13], X[13], Y[13]);
  GPGenerator U5 (G0[14], P0[14], X[14], Y[14]);
  GPGenerator U6 (G0[15], P0[15], X[15], Y[15]);
  GPGenerator U7 (G0[16], P0[16], X[16], Y[16]);
  GPGenerator U8 (G0[17], P0[17], X[17], Y[17]);
  GPGenerator U9 (G0[18], P0[18], X[18], Y[18]);
  GPGenerator U10 (G0[19], P0[19], X[19], Y[19]);
  GPGenerator U11 (G0[20], P0[20], X[20], Y[20]);
  GPGenerator U12 (G0[21], P0[21], X[21], Y[21]);
  GPGenerator U13 (G0[22], P0[22], X[22], Y[22]);
  GPGenerator U14 (G0[23], P0[23], X[23], Y[23]);
  GPGenerator U15 (G0[24], P0[24], X[24], Y[24]);
  GPGenerator U16 (G0[25], P0[25], X[25], Y[25]);
  GPGenerator U17 (G0[26], P0[26], X[26], Y[26]);
  GPGenerator U18 (G0[27], P0[27], X[27], Y[27]);
  GPGenerator U19 (G0[28], P0[28], X[28], Y[28]);
  GPGenerator U20 (G0[29], P0[29], X[29], Y[29]);
  GPGenerator U21 (G0[30], P0[30], X[30], Y[30]);
  GPGenerator U22 (G0[31], P0[31], X[31], Y[31]);
  GPGenerator U23 (G0[32], P0[32], X[32], Y[32]);
  GPGenerator U24 (G0[33], P0[33], X[33], Y[33]);
  GPGenerator U25 (G0[34], P0[34], X[34], Y[34]);
  GPGenerator U26 (G0[35], P0[35], X[35], Y[35]);
  GPGenerator U27 (G0[36], P0[36], X[36], Y[36]);
  GPGenerator U28 (G0[37], P0[37], X[37], Y[37]);
  GPGenerator U29 (G0[38], P0[38], X[38], Y[38]);
  GPGenerator U30 (G0[39], P0[39], X[39], Y[39]);
  GPGenerator U31 (G0[40], P0[40], X[40], Y[40]);
  GPGenerator U32 (G0[41], P0[41], X[41], Y[41]);
  GPGenerator U33 (G0[42], P0[42], X[42], Y[42]);
  GPGenerator U34 (G0[43], P0[43], X[43], Y[43]);
  GPGenerator U35 (G0[44], P0[44], X[44], Y[44]);
  GPGenerator U36 (G0[45], P0[45], X[45], Y[45]);
  GPGenerator U37 (G0[46], P0[46], X[46], Y[46]);
  GPGenerator U38 (G0[47], P0[47], X[47], Y[47]);
  GPGenerator U39 (G0[48], P0[48], X[48], Y[48]);
  GPGenerator U40 (G0[49], P0[49], X[49], Y[49]);
  GPGenerator U41 (G0[50], P0[50], X[50], Y[50]);
  GPGenerator U42 (G0[51], P0[51], X[51], Y[51]);
  GPGenerator U43 (G0[52], P0[52], X[52], Y[52]);
  GPGenerator U44 (G0[53], P0[53], X[53], Y[53]);
  GPGenerator U45 (G0[54], P0[54], X[54], Y[54]);
  GPGenerator U46 (G0[55], P0[55], X[55], Y[55]);
  GPGenerator U47 (G0[56], P0[56], X[56], Y[56]);
  GPGenerator U48 (G0[57], P0[57], X[57], Y[57]);
  GPGenerator U49 (G0[58], P0[58], X[58], Y[58]);
  GPGenerator U50 (G0[59], P0[59], X[59], Y[59]);
  GPGenerator U51 (G0[60], P0[60], X[60], Y[60]);
  GPGenerator U52 (G0[61], P0[61], X[61], Y[61]);
  GPGenerator U53 (G0[62], P0[62], X[62], Y[62]);
  GPGenerator U54 (G0[63], P0[63], X[63], Y[63]);
  GPGenerator U55 (G0[64], P0[64], X[64], Y[64]);
  CarryOperator U56 (G1[10], P1[10], G0[10], P0[10], G0[9], P0[9]);
  CarryOperator U57 (G1[11], P1[11], G0[11], P0[11], G0[10], P0[10]);
  CarryOperator U58 (G1[12], P1[12], G0[12], P0[12], G0[11], P0[11]);
  CarryOperator U59 (G1[13], P1[13], G0[13], P0[13], G0[12], P0[12]);
  CarryOperator U60 (G1[14], P1[14], G0[14], P0[14], G0[13], P0[13]);
  CarryOperator U61 (G1[15], P1[15], G0[15], P0[15], G0[14], P0[14]);
  CarryOperator U62 (G1[16], P1[16], G0[16], P0[16], G0[15], P0[15]);
  CarryOperator U63 (G1[17], P1[17], G0[17], P0[17], G0[16], P0[16]);
  CarryOperator U64 (G1[18], P1[18], G0[18], P0[18], G0[17], P0[17]);
  CarryOperator U65 (G1[19], P1[19], G0[19], P0[19], G0[18], P0[18]);
  CarryOperator U66 (G1[20], P1[20], G0[20], P0[20], G0[19], P0[19]);
  CarryOperator U67 (G1[21], P1[21], G0[21], P0[21], G0[20], P0[20]);
  CarryOperator U68 (G1[22], P1[22], G0[22], P0[22], G0[21], P0[21]);
  CarryOperator U69 (G1[23], P1[23], G0[23], P0[23], G0[22], P0[22]);
  CarryOperator U70 (G1[24], P1[24], G0[24], P0[24], G0[23], P0[23]);
  CarryOperator U71 (G1[25], P1[25], G0[25], P0[25], G0[24], P0[24]);
  CarryOperator U72 (G1[26], P1[26], G0[26], P0[26], G0[25], P0[25]);
  CarryOperator U73 (G1[27], P1[27], G0[27], P0[27], G0[26], P0[26]);
  CarryOperator U74 (G1[28], P1[28], G0[28], P0[28], G0[27], P0[27]);
  CarryOperator U75 (G1[29], P1[29], G0[29], P0[29], G0[28], P0[28]);
  CarryOperator U76 (G1[30], P1[30], G0[30], P0[30], G0[29], P0[29]);
  CarryOperator U77 (G1[31], P1[31], G0[31], P0[31], G0[30], P0[30]);
  CarryOperator U78 (G1[32], P1[32], G0[32], P0[32], G0[31], P0[31]);
  CarryOperator U79 (G1[33], P1[33], G0[33], P0[33], G0[32], P0[32]);
  CarryOperator U80 (G1[34], P1[34], G0[34], P0[34], G0[33], P0[33]);
  CarryOperator U81 (G1[35], P1[35], G0[35], P0[35], G0[34], P0[34]);
  CarryOperator U82 (G1[36], P1[36], G0[36], P0[36], G0[35], P0[35]);
  CarryOperator U83 (G1[37], P1[37], G0[37], P0[37], G0[36], P0[36]);
  CarryOperator U84 (G1[38], P1[38], G0[38], P0[38], G0[37], P0[37]);
  CarryOperator U85 (G1[39], P1[39], G0[39], P0[39], G0[38], P0[38]);
  CarryOperator U86 (G1[40], P1[40], G0[40], P0[40], G0[39], P0[39]);
  CarryOperator U87 (G1[41], P1[41], G0[41], P0[41], G0[40], P0[40]);
  CarryOperator U88 (G1[42], P1[42], G0[42], P0[42], G0[41], P0[41]);
  CarryOperator U89 (G1[43], P1[43], G0[43], P0[43], G0[42], P0[42]);
  CarryOperator U90 (G1[44], P1[44], G0[44], P0[44], G0[43], P0[43]);
  CarryOperator U91 (G1[45], P1[45], G0[45], P0[45], G0[44], P0[44]);
  CarryOperator U92 (G1[46], P1[46], G0[46], P0[46], G0[45], P0[45]);
  CarryOperator U93 (G1[47], P1[47], G0[47], P0[47], G0[46], P0[46]);
  CarryOperator U94 (G1[48], P1[48], G0[48], P0[48], G0[47], P0[47]);
  CarryOperator U95 (G1[49], P1[49], G0[49], P0[49], G0[48], P0[48]);
  CarryOperator U96 (G1[50], P1[50], G0[50], P0[50], G0[49], P0[49]);
  CarryOperator U97 (G1[51], P1[51], G0[51], P0[51], G0[50], P0[50]);
  CarryOperator U98 (G1[52], P1[52], G0[52], P0[52], G0[51], P0[51]);
  CarryOperator U99 (G1[53], P1[53], G0[53], P0[53], G0[52], P0[52]);
  CarryOperator U100 (G1[54], P1[54], G0[54], P0[54], G0[53], P0[53]);
  CarryOperator U101 (G1[55], P1[55], G0[55], P0[55], G0[54], P0[54]);
  CarryOperator U102 (G1[56], P1[56], G0[56], P0[56], G0[55], P0[55]);
  CarryOperator U103 (G1[57], P1[57], G0[57], P0[57], G0[56], P0[56]);
  CarryOperator U104 (G1[58], P1[58], G0[58], P0[58], G0[57], P0[57]);
  CarryOperator U105 (G1[59], P1[59], G0[59], P0[59], G0[58], P0[58]);
  CarryOperator U106 (G1[60], P1[60], G0[60], P0[60], G0[59], P0[59]);
  CarryOperator U107 (G1[61], P1[61], G0[61], P0[61], G0[60], P0[60]);
  CarryOperator U108 (G1[62], P1[62], G0[62], P0[62], G0[61], P0[61]);
  CarryOperator U109 (G1[63], P1[63], G0[63], P0[63], G0[62], P0[62]);
  CarryOperator U110 (G1[64], P1[64], G0[64], P0[64], G0[63], P0[63]);
  CarryOperator U111 (G2[11], P2[11], G1[11], P1[11], G1[9], P1[9]);
  CarryOperator U112 (G2[12], P2[12], G1[12], P1[12], G1[10], P1[10]);
  CarryOperator U113 (G2[13], P2[13], G1[13], P1[13], G1[11], P1[11]);
  CarryOperator U114 (G2[14], P2[14], G1[14], P1[14], G1[12], P1[12]);
  CarryOperator U115 (G2[15], P2[15], G1[15], P1[15], G1[13], P1[13]);
  CarryOperator U116 (G2[16], P2[16], G1[16], P1[16], G1[14], P1[14]);
  CarryOperator U117 (G2[17], P2[17], G1[17], P1[17], G1[15], P1[15]);
  CarryOperator U118 (G2[18], P2[18], G1[18], P1[18], G1[16], P1[16]);
  CarryOperator U119 (G2[19], P2[19], G1[19], P1[19], G1[17], P1[17]);
  CarryOperator U120 (G2[20], P2[20], G1[20], P1[20], G1[18], P1[18]);
  CarryOperator U121 (G2[21], P2[21], G1[21], P1[21], G1[19], P1[19]);
  CarryOperator U122 (G2[22], P2[22], G1[22], P1[22], G1[20], P1[20]);
  CarryOperator U123 (G2[23], P2[23], G1[23], P1[23], G1[21], P1[21]);
  CarryOperator U124 (G2[24], P2[24], G1[24], P1[24], G1[22], P1[22]);
  CarryOperator U125 (G2[25], P2[25], G1[25], P1[25], G1[23], P1[23]);
  CarryOperator U126 (G2[26], P2[26], G1[26], P1[26], G1[24], P1[24]);
  CarryOperator U127 (G2[27], P2[27], G1[27], P1[27], G1[25], P1[25]);
  CarryOperator U128 (G2[28], P2[28], G1[28], P1[28], G1[26], P1[26]);
  CarryOperator U129 (G2[29], P2[29], G1[29], P1[29], G1[27], P1[27]);
  CarryOperator U130 (G2[30], P2[30], G1[30], P1[30], G1[28], P1[28]);
  CarryOperator U131 (G2[31], P2[31], G1[31], P1[31], G1[29], P1[29]);
  CarryOperator U132 (G2[32], P2[32], G1[32], P1[32], G1[30], P1[30]);
  CarryOperator U133 (G2[33], P2[33], G1[33], P1[33], G1[31], P1[31]);
  CarryOperator U134 (G2[34], P2[34], G1[34], P1[34], G1[32], P1[32]);
  CarryOperator U135 (G2[35], P2[35], G1[35], P1[35], G1[33], P1[33]);
  CarryOperator U136 (G2[36], P2[36], G1[36], P1[36], G1[34], P1[34]);
  CarryOperator U137 (G2[37], P2[37], G1[37], P1[37], G1[35], P1[35]);
  CarryOperator U138 (G2[38], P2[38], G1[38], P1[38], G1[36], P1[36]);
  CarryOperator U139 (G2[39], P2[39], G1[39], P1[39], G1[37], P1[37]);
  CarryOperator U140 (G2[40], P2[40], G1[40], P1[40], G1[38], P1[38]);
  CarryOperator U141 (G2[41], P2[41], G1[41], P1[41], G1[39], P1[39]);
  CarryOperator U142 (G2[42], P2[42], G1[42], P1[42], G1[40], P1[40]);
  CarryOperator U143 (G2[43], P2[43], G1[43], P1[43], G1[41], P1[41]);
  CarryOperator U144 (G2[44], P2[44], G1[44], P1[44], G1[42], P1[42]);
  CarryOperator U145 (G2[45], P2[45], G1[45], P1[45], G1[43], P1[43]);
  CarryOperator U146 (G2[46], P2[46], G1[46], P1[46], G1[44], P1[44]);
  CarryOperator U147 (G2[47], P2[47], G1[47], P1[47], G1[45], P1[45]);
  CarryOperator U148 (G2[48], P2[48], G1[48], P1[48], G1[46], P1[46]);
  CarryOperator U149 (G2[49], P2[49], G1[49], P1[49], G1[47], P1[47]);
  CarryOperator U150 (G2[50], P2[50], G1[50], P1[50], G1[48], P1[48]);
  CarryOperator U151 (G2[51], P2[51], G1[51], P1[51], G1[49], P1[49]);
  CarryOperator U152 (G2[52], P2[52], G1[52], P1[52], G1[50], P1[50]);
  CarryOperator U153 (G2[53], P2[53], G1[53], P1[53], G1[51], P1[51]);
  CarryOperator U154 (G2[54], P2[54], G1[54], P1[54], G1[52], P1[52]);
  CarryOperator U155 (G2[55], P2[55], G1[55], P1[55], G1[53], P1[53]);
  CarryOperator U156 (G2[56], P2[56], G1[56], P1[56], G1[54], P1[54]);
  CarryOperator U157 (G2[57], P2[57], G1[57], P1[57], G1[55], P1[55]);
  CarryOperator U158 (G2[58], P2[58], G1[58], P1[58], G1[56], P1[56]);
  CarryOperator U159 (G2[59], P2[59], G1[59], P1[59], G1[57], P1[57]);
  CarryOperator U160 (G2[60], P2[60], G1[60], P1[60], G1[58], P1[58]);
  CarryOperator U161 (G2[61], P2[61], G1[61], P1[61], G1[59], P1[59]);
  CarryOperator U162 (G2[62], P2[62], G1[62], P1[62], G1[60], P1[60]);
  CarryOperator U163 (G2[63], P2[63], G1[63], P1[63], G1[61], P1[61]);
  CarryOperator U164 (G2[64], P2[64], G1[64], P1[64], G1[62], P1[62]);
  CarryOperator U165 (G3[13], P3[13], G2[13], P2[13], G2[9], P2[9]);
  CarryOperator U166 (G3[14], P3[14], G2[14], P2[14], G2[10], P2[10]);
  CarryOperator U167 (G3[15], P3[15], G2[15], P2[15], G2[11], P2[11]);
  CarryOperator U168 (G3[16], P3[16], G2[16], P2[16], G2[12], P2[12]);
  CarryOperator U169 (G3[17], P3[17], G2[17], P2[17], G2[13], P2[13]);
  CarryOperator U170 (G3[18], P3[18], G2[18], P2[18], G2[14], P2[14]);
  CarryOperator U171 (G3[19], P3[19], G2[19], P2[19], G2[15], P2[15]);
  CarryOperator U172 (G3[20], P3[20], G2[20], P2[20], G2[16], P2[16]);
  CarryOperator U173 (G3[21], P3[21], G2[21], P2[21], G2[17], P2[17]);
  CarryOperator U174 (G3[22], P3[22], G2[22], P2[22], G2[18], P2[18]);
  CarryOperator U175 (G3[23], P3[23], G2[23], P2[23], G2[19], P2[19]);
  CarryOperator U176 (G3[24], P3[24], G2[24], P2[24], G2[20], P2[20]);
  CarryOperator U177 (G3[25], P3[25], G2[25], P2[25], G2[21], P2[21]);
  CarryOperator U178 (G3[26], P3[26], G2[26], P2[26], G2[22], P2[22]);
  CarryOperator U179 (G3[27], P3[27], G2[27], P2[27], G2[23], P2[23]);
  CarryOperator U180 (G3[28], P3[28], G2[28], P2[28], G2[24], P2[24]);
  CarryOperator U181 (G3[29], P3[29], G2[29], P2[29], G2[25], P2[25]);
  CarryOperator U182 (G3[30], P3[30], G2[30], P2[30], G2[26], P2[26]);
  CarryOperator U183 (G3[31], P3[31], G2[31], P2[31], G2[27], P2[27]);
  CarryOperator U184 (G3[32], P3[32], G2[32], P2[32], G2[28], P2[28]);
  CarryOperator U185 (G3[33], P3[33], G2[33], P2[33], G2[29], P2[29]);
  CarryOperator U186 (G3[34], P3[34], G2[34], P2[34], G2[30], P2[30]);
  CarryOperator U187 (G3[35], P3[35], G2[35], P2[35], G2[31], P2[31]);
  CarryOperator U188 (G3[36], P3[36], G2[36], P2[36], G2[32], P2[32]);
  CarryOperator U189 (G3[37], P3[37], G2[37], P2[37], G2[33], P2[33]);
  CarryOperator U190 (G3[38], P3[38], G2[38], P2[38], G2[34], P2[34]);
  CarryOperator U191 (G3[39], P3[39], G2[39], P2[39], G2[35], P2[35]);
  CarryOperator U192 (G3[40], P3[40], G2[40], P2[40], G2[36], P2[36]);
  CarryOperator U193 (G3[41], P3[41], G2[41], P2[41], G2[37], P2[37]);
  CarryOperator U194 (G3[42], P3[42], G2[42], P2[42], G2[38], P2[38]);
  CarryOperator U195 (G3[43], P3[43], G2[43], P2[43], G2[39], P2[39]);
  CarryOperator U196 (G3[44], P3[44], G2[44], P2[44], G2[40], P2[40]);
  CarryOperator U197 (G3[45], P3[45], G2[45], P2[45], G2[41], P2[41]);
  CarryOperator U198 (G3[46], P3[46], G2[46], P2[46], G2[42], P2[42]);
  CarryOperator U199 (G3[47], P3[47], G2[47], P2[47], G2[43], P2[43]);
  CarryOperator U200 (G3[48], P3[48], G2[48], P2[48], G2[44], P2[44]);
  CarryOperator U201 (G3[49], P3[49], G2[49], P2[49], G2[45], P2[45]);
  CarryOperator U202 (G3[50], P3[50], G2[50], P2[50], G2[46], P2[46]);
  CarryOperator U203 (G3[51], P3[51], G2[51], P2[51], G2[47], P2[47]);
  CarryOperator U204 (G3[52], P3[52], G2[52], P2[52], G2[48], P2[48]);
  CarryOperator U205 (G3[53], P3[53], G2[53], P2[53], G2[49], P2[49]);
  CarryOperator U206 (G3[54], P3[54], G2[54], P2[54], G2[50], P2[50]);
  CarryOperator U207 (G3[55], P3[55], G2[55], P2[55], G2[51], P2[51]);
  CarryOperator U208 (G3[56], P3[56], G2[56], P2[56], G2[52], P2[52]);
  CarryOperator U209 (G3[57], P3[57], G2[57], P2[57], G2[53], P2[53]);
  CarryOperator U210 (G3[58], P3[58], G2[58], P2[58], G2[54], P2[54]);
  CarryOperator U211 (G3[59], P3[59], G2[59], P2[59], G2[55], P2[55]);
  CarryOperator U212 (G3[60], P3[60], G2[60], P2[60], G2[56], P2[56]);
  CarryOperator U213 (G3[61], P3[61], G2[61], P2[61], G2[57], P2[57]);
  CarryOperator U214 (G3[62], P3[62], G2[62], P2[62], G2[58], P2[58]);
  CarryOperator U215 (G3[63], P3[63], G2[63], P2[63], G2[59], P2[59]);
  CarryOperator U216 (G3[64], P3[64], G2[64], P2[64], G2[60], P2[60]);
  CarryOperator U217 (G4[17], P4[17], G3[17], P3[17], G3[9], P3[9]);
  CarryOperator U218 (G4[18], P4[18], G3[18], P3[18], G3[10], P3[10]);
  CarryOperator U219 (G4[19], P4[19], G3[19], P3[19], G3[11], P3[11]);
  CarryOperator U220 (G4[20], P4[20], G3[20], P3[20], G3[12], P3[12]);
  CarryOperator U221 (G4[21], P4[21], G3[21], P3[21], G3[13], P3[13]);
  CarryOperator U222 (G4[22], P4[22], G3[22], P3[22], G3[14], P3[14]);
  CarryOperator U223 (G4[23], P4[23], G3[23], P3[23], G3[15], P3[15]);
  CarryOperator U224 (G4[24], P4[24], G3[24], P3[24], G3[16], P3[16]);
  CarryOperator U225 (G4[25], P4[25], G3[25], P3[25], G3[17], P3[17]);
  CarryOperator U226 (G4[26], P4[26], G3[26], P3[26], G3[18], P3[18]);
  CarryOperator U227 (G4[27], P4[27], G3[27], P3[27], G3[19], P3[19]);
  CarryOperator U228 (G4[28], P4[28], G3[28], P3[28], G3[20], P3[20]);
  CarryOperator U229 (G4[29], P4[29], G3[29], P3[29], G3[21], P3[21]);
  CarryOperator U230 (G4[30], P4[30], G3[30], P3[30], G3[22], P3[22]);
  CarryOperator U231 (G4[31], P4[31], G3[31], P3[31], G3[23], P3[23]);
  CarryOperator U232 (G4[32], P4[32], G3[32], P3[32], G3[24], P3[24]);
  CarryOperator U233 (G4[33], P4[33], G3[33], P3[33], G3[25], P3[25]);
  CarryOperator U234 (G4[34], P4[34], G3[34], P3[34], G3[26], P3[26]);
  CarryOperator U235 (G4[35], P4[35], G3[35], P3[35], G3[27], P3[27]);
  CarryOperator U236 (G4[36], P4[36], G3[36], P3[36], G3[28], P3[28]);
  CarryOperator U237 (G4[37], P4[37], G3[37], P3[37], G3[29], P3[29]);
  CarryOperator U238 (G4[38], P4[38], G3[38], P3[38], G3[30], P3[30]);
  CarryOperator U239 (G4[39], P4[39], G3[39], P3[39], G3[31], P3[31]);
  CarryOperator U240 (G4[40], P4[40], G3[40], P3[40], G3[32], P3[32]);
  CarryOperator U241 (G4[41], P4[41], G3[41], P3[41], G3[33], P3[33]);
  CarryOperator U242 (G4[42], P4[42], G3[42], P3[42], G3[34], P3[34]);
  CarryOperator U243 (G4[43], P4[43], G3[43], P3[43], G3[35], P3[35]);
  CarryOperator U244 (G4[44], P4[44], G3[44], P3[44], G3[36], P3[36]);
  CarryOperator U245 (G4[45], P4[45], G3[45], P3[45], G3[37], P3[37]);
  CarryOperator U246 (G4[46], P4[46], G3[46], P3[46], G3[38], P3[38]);
  CarryOperator U247 (G4[47], P4[47], G3[47], P3[47], G3[39], P3[39]);
  CarryOperator U248 (G4[48], P4[48], G3[48], P3[48], G3[40], P3[40]);
  CarryOperator U249 (G4[49], P4[49], G3[49], P3[49], G3[41], P3[41]);
  CarryOperator U250 (G4[50], P4[50], G3[50], P3[50], G3[42], P3[42]);
  CarryOperator U251 (G4[51], P4[51], G3[51], P3[51], G3[43], P3[43]);
  CarryOperator U252 (G4[52], P4[52], G3[52], P3[52], G3[44], P3[44]);
  CarryOperator U253 (G4[53], P4[53], G3[53], P3[53], G3[45], P3[45]);
  CarryOperator U254 (G4[54], P4[54], G3[54], P3[54], G3[46], P3[46]);
  CarryOperator U255 (G4[55], P4[55], G3[55], P3[55], G3[47], P3[47]);
  CarryOperator U256 (G4[56], P4[56], G3[56], P3[56], G3[48], P3[48]);
  CarryOperator U257 (G4[57], P4[57], G3[57], P3[57], G3[49], P3[49]);
  CarryOperator U258 (G4[58], P4[58], G3[58], P3[58], G3[50], P3[50]);
  CarryOperator U259 (G4[59], P4[59], G3[59], P3[59], G3[51], P3[51]);
  CarryOperator U260 (G4[60], P4[60], G3[60], P3[60], G3[52], P3[52]);
  CarryOperator U261 (G4[61], P4[61], G3[61], P3[61], G3[53], P3[53]);
  CarryOperator U262 (G4[62], P4[62], G3[62], P3[62], G3[54], P3[54]);
  CarryOperator U263 (G4[63], P4[63], G3[63], P3[63], G3[55], P3[55]);
  CarryOperator U264 (G4[64], P4[64], G3[64], P3[64], G3[56], P3[56]);
  CarryOperator U265 (G5[25], P5[25], G4[25], P4[25], G4[9], P4[9]);
  CarryOperator U266 (G5[26], P5[26], G4[26], P4[26], G4[10], P4[10]);
  CarryOperator U267 (G5[27], P5[27], G4[27], P4[27], G4[11], P4[11]);
  CarryOperator U268 (G5[28], P5[28], G4[28], P4[28], G4[12], P4[12]);
  CarryOperator U269 (G5[29], P5[29], G4[29], P4[29], G4[13], P4[13]);
  CarryOperator U270 (G5[30], P5[30], G4[30], P4[30], G4[14], P4[14]);
  CarryOperator U271 (G5[31], P5[31], G4[31], P4[31], G4[15], P4[15]);
  CarryOperator U272 (G5[32], P5[32], G4[32], P4[32], G4[16], P4[16]);
  CarryOperator U273 (G5[33], P5[33], G4[33], P4[33], G4[17], P4[17]);
  CarryOperator U274 (G5[34], P5[34], G4[34], P4[34], G4[18], P4[18]);
  CarryOperator U275 (G5[35], P5[35], G4[35], P4[35], G4[19], P4[19]);
  CarryOperator U276 (G5[36], P5[36], G4[36], P4[36], G4[20], P4[20]);
  CarryOperator U277 (G5[37], P5[37], G4[37], P4[37], G4[21], P4[21]);
  CarryOperator U278 (G5[38], P5[38], G4[38], P4[38], G4[22], P4[22]);
  CarryOperator U279 (G5[39], P5[39], G4[39], P4[39], G4[23], P4[23]);
  CarryOperator U280 (G5[40], P5[40], G4[40], P4[40], G4[24], P4[24]);
  CarryOperator U281 (G5[41], P5[41], G4[41], P4[41], G4[25], P4[25]);
  CarryOperator U282 (G5[42], P5[42], G4[42], P4[42], G4[26], P4[26]);
  CarryOperator U283 (G5[43], P5[43], G4[43], P4[43], G4[27], P4[27]);
  CarryOperator U284 (G5[44], P5[44], G4[44], P4[44], G4[28], P4[28]);
  CarryOperator U285 (G5[45], P5[45], G4[45], P4[45], G4[29], P4[29]);
  CarryOperator U286 (G5[46], P5[46], G4[46], P4[46], G4[30], P4[30]);
  CarryOperator U287 (G5[47], P5[47], G4[47], P4[47], G4[31], P4[31]);
  CarryOperator U288 (G5[48], P5[48], G4[48], P4[48], G4[32], P4[32]);
  CarryOperator U289 (G5[49], P5[49], G4[49], P4[49], G4[33], P4[33]);
  CarryOperator U290 (G5[50], P5[50], G4[50], P4[50], G4[34], P4[34]);
  CarryOperator U291 (G5[51], P5[51], G4[51], P4[51], G4[35], P4[35]);
  CarryOperator U292 (G5[52], P5[52], G4[52], P4[52], G4[36], P4[36]);
  CarryOperator U293 (G5[53], P5[53], G4[53], P4[53], G4[37], P4[37]);
  CarryOperator U294 (G5[54], P5[54], G4[54], P4[54], G4[38], P4[38]);
  CarryOperator U295 (G5[55], P5[55], G4[55], P4[55], G4[39], P4[39]);
  CarryOperator U296 (G5[56], P5[56], G4[56], P4[56], G4[40], P4[40]);
  CarryOperator U297 (G5[57], P5[57], G4[57], P4[57], G4[41], P4[41]);
  CarryOperator U298 (G5[58], P5[58], G4[58], P4[58], G4[42], P4[42]);
  CarryOperator U299 (G5[59], P5[59], G4[59], P4[59], G4[43], P4[43]);
  CarryOperator U300 (G5[60], P5[60], G4[60], P4[60], G4[44], P4[44]);
  CarryOperator U301 (G5[61], P5[61], G4[61], P4[61], G4[45], P4[45]);
  CarryOperator U302 (G5[62], P5[62], G4[62], P4[62], G4[46], P4[46]);
  CarryOperator U303 (G5[63], P5[63], G4[63], P4[63], G4[47], P4[47]);
  CarryOperator U304 (G5[64], P5[64], G4[64], P4[64], G4[48], P4[48]);
  CarryOperator U305 (G6[41], P6[41], G5[41], P5[41], G5[9], P5[9]);
  CarryOperator U306 (G6[42], P6[42], G5[42], P5[42], G5[10], P5[10]);
  CarryOperator U307 (G6[43], P6[43], G5[43], P5[43], G5[11], P5[11]);
  CarryOperator U308 (G6[44], P6[44], G5[44], P5[44], G5[12], P5[12]);
  CarryOperator U309 (G6[45], P6[45], G5[45], P5[45], G5[13], P5[13]);
  CarryOperator U310 (G6[46], P6[46], G5[46], P5[46], G5[14], P5[14]);
  CarryOperator U311 (G6[47], P6[47], G5[47], P5[47], G5[15], P5[15]);
  CarryOperator U312 (G6[48], P6[48], G5[48], P5[48], G5[16], P5[16]);
  CarryOperator U313 (G6[49], P6[49], G5[49], P5[49], G5[17], P5[17]);
  CarryOperator U314 (G6[50], P6[50], G5[50], P5[50], G5[18], P5[18]);
  CarryOperator U315 (G6[51], P6[51], G5[51], P5[51], G5[19], P5[19]);
  CarryOperator U316 (G6[52], P6[52], G5[52], P5[52], G5[20], P5[20]);
  CarryOperator U317 (G6[53], P6[53], G5[53], P5[53], G5[21], P5[21]);
  CarryOperator U318 (G6[54], P6[54], G5[54], P5[54], G5[22], P5[22]);
  CarryOperator U319 (G6[55], P6[55], G5[55], P5[55], G5[23], P5[23]);
  CarryOperator U320 (G6[56], P6[56], G5[56], P5[56], G5[24], P5[24]);
  CarryOperator U321 (G6[57], P6[57], G5[57], P5[57], G5[25], P5[25]);
  CarryOperator U322 (G6[58], P6[58], G5[58], P5[58], G5[26], P5[26]);
  CarryOperator U323 (G6[59], P6[59], G5[59], P5[59], G5[27], P5[27]);
  CarryOperator U324 (G6[60], P6[60], G5[60], P5[60], G5[28], P5[28]);
  CarryOperator U325 (G6[61], P6[61], G5[61], P5[61], G5[29], P5[29]);
  CarryOperator U326 (G6[62], P6[62], G5[62], P5[62], G5[30], P5[30]);
  CarryOperator U327 (G6[63], P6[63], G5[63], P5[63], G5[31], P5[31]);
  CarryOperator U328 (G6[64], P6[64], G5[64], P5[64], G5[32], P5[32]);
endmodule

module UBZero_9_9(O);
  output [9:9] O;
  assign O[9] = 0;
endmodule

module UBTC1CON66_0(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_1(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_2(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_3(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_4(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_5(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_6(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_7(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_8(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_9(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_10(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_11(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_12(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_13(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_14(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_15(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_16(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_17(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_18(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_19(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_20(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_21(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_22(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_23(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_24(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_25(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_26(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_27(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_28(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_29(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_30(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_31(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_32(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_33(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_34(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_35(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_36(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_37(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_38(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_39(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_40(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_41(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_42(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_43(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_44(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_45(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_46(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_47(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_48(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_49(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_50(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_51(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_52(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_53(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_54(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_55(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_56(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_57(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_58(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_59(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_60(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_61(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTC1CON66_62(O, I);
  output O;
  input I;
  assign O = I;
endmodule

module UBTCTCONV_65_63(O, I);
  output [66:63] O;
  input [65:63] I;
  assign O[63] = ~ I[63];
  assign O[64] = ~ I[64] ^ ( I[63] );
  assign O[65] = ~ I[65] ^ ( I[64] | I[63] );
  assign O[66] = ~ ( I[65] | I[64] | I[63] );
endmodule

module multiplier_32b(P, IN1, IN2, clk, rst);

  input clk, rst;
  
  output [63:0] P;
  reg [63:0] P_reg;
  input [31:0] IN1;
  input [31:0] IN2;
  wire [66:0] W;

  reg [31:0]  IN1_reg;
  reg [31:0]  IN2_reg;
   
  always @(posedge clk)
  begin
		if(rst)
		begin
			IN1_reg <= 0;
			IN2_reg <= 0;
			P_reg 	<= 0;
		end
		else
		begin
			IN1_reg <= IN1;
			IN2_reg <= IN2;
			P_reg   <= W[63:0];
		end
  end
   
  assign P = P_reg; 
   

  //assign P[0] = W[0];
  //assign P[1] = W[1];
  //assign P[2] = W[2];
  //assign P[3] = W[3];
  //assign P[4] = W[4];
  //assign P[5] = W[5];
  //assign P[6] = W[6];
  //assign P[7] = W[7];
  //assign P[8] = W[8];
  //assign P[9] = W[9];
  //assign P[10] = W[10];
  //assign P[11] = W[11];
  //assign P[12] = W[12];
  //assign P[13] = W[13];
  //assign P[14] = W[14];
  //assign P[15] = W[15];
  //assign P[16] = W[16];
  //assign P[17] = W[17];
  //assign P[18] = W[18];
  //assign P[19] = W[19];
  //assign P[20] = W[20];
  //assign P[21] = W[21];
  //assign P[22] = W[22];
  //assign P[23] = W[23];
  //assign P[24] = W[24];
  //assign P[25] = W[25];
  //assign P[26] = W[26];
  //assign P[27] = W[27];
  //assign P[28] = W[28];
  //assign P[29] = W[29];
  //assign P[30] = W[30];
  //assign P[31] = W[31];
  //assign P[32] = W[32];
  //assign P[33] = W[33];
  //assign P[34] = W[34];
  //assign P[35] = W[35];
  //assign P[36] = W[36];
  //assign P[37] = W[37];
  //assign P[38] = W[38];
  //assign P[39] = W[39];
  //assign P[40] = W[40];
  //assign P[41] = W[41];
  //assign P[42] = W[42];
  //assign P[43] = W[43];
  //assign P[44] = W[44];
  //assign P[45] = W[45];
  //assign P[46] = W[46];
  //assign P[47] = W[47];
  //assign P[48] = W[48];
  //assign P[49] = W[49];
  //assign P[50] = W[50];
  //assign P[51] = W[51];
  //assign P[52] = W[52];
  //assign P[53] = W[53];
  //assign P[54] = W[54];
  //assign P[55] = W[55];
  //assign P[56] = W[56];
  //assign P[57] = W[57];
  //assign P[58] = W[58];
  //assign P[59] = W[59];
  //assign P[60] = W[60];
  //assign P[61] = W[61];
  //assign P[62] = W[62];
  //assign P[63] = W[63];

  MultTC_STD_WAL_KS000 U0 (W, IN1_reg, IN2_reg, clk, rst);
endmodule

module CSA_32_0_32_1_33_000 (C, S, X, Y, Z);
  output [33:2] C;
  output [33:0] S;
  input [32:0] X;
  input [32:1] Y;
  input [33:2] Z;
  UB1DCON_0 U0 (S[0], X[0]);
  UBHA_1 U1 (C[2], S[1], Y[1], X[1]);
  PureCSA_32_2 U2 (C[33:3], S[32:2], Z[32:2], Y[32:2], X[32:2]);
  UB1DCON_33 U3 (S[33], Z[33]);
endmodule

module CSA_33_0_33_2_36_000 (C, S, X, Y, Z);
  output [34:3] C;
  output [36:0] S;
  input [33:0] X;
  input [33:2] Y;
  input [36:3] Z;
  UBCON_1_0 U0 (S[1:0], X[1:0]);
  UBHA_2 U1 (C[3], S[2], Y[2], X[2]);
  PureCSA_33_3 U2 (C[34:4], S[33:3], Z[33:3], Y[33:3], X[33:3]);
  UBCON_36_34 U3 (S[36:34], Z[36:34]);
endmodule

module CSA_34_3_35_4_36_000 (C, S, X, Y, Z);
  output [36:5] C;
  output [36:3] S;
  input [34:3] X;
  input [35:4] Y;
  input [36:5] Z;
  UB1DCON_3 U0 (S[3], X[3]);
  UBHA_4 U1 (C[5], S[4], Y[4], X[4]);
  PureCSA_34_5 U2 (C[35:6], S[34:5], Z[34:5], Y[34:5], X[34:5]);
  UBHA_35 U3 (C[36], S[35], Z[35], Y[35]);
  UB1DCON_36 U4 (S[36], Z[36]);
endmodule

module CSA_36_0_34_3_39_000 (C, S, X, Y, Z);
  output [37:4] C;
  output [39:0] S;
  input [36:0] X;
  input [34:3] Y;
  input [39:5] Z;
  UBCON_2_0 U0 (S[2:0], X[2:0]);
  PureCSHA_4_3 U1 (C[5:4], S[4:3], Y[4:3], X[4:3]);
  PureCSA_34_5 U2 (C[35:6], S[34:5], Z[34:5], Y[34:5], X[34:5]);
  PureCSHA_36_35 U3 (C[37:36], S[36:35], Z[36:35], X[36:35]);
  UBCON_39_37 U4 (S[39:37], Z[39:37]);
endmodule

module CSA_36_5_39_6_39_000 (C, S, X, Y, Z);
  output [40:7] C;
  output [39:5] S;
  input [36:5] X;
  input [39:6] Y;
  input [39:8] Z;
  UB1DCON_5 U0 (S[5], X[5]);
  PureCSHA_7_6 U1 (C[8:7], S[7:6], Y[7:6], X[7:6]);
  PureCSA_36_8 U2 (C[37:9], S[36:8], Z[36:8], Y[36:8], X[36:8]);
  PureCSHA_39_37 U3 (C[40:38], S[39:37], Z[39:37], Y[39:37]);
endmodule

module CSA_37_6_38_7_39_000 (C, S, X, Y, Z);
  output [39:8] C;
  output [39:6] S;
  input [37:6] X;
  input [38:7] Y;
  input [39:8] Z;
  UB1DCON_6 U0 (S[6], X[6]);
  UBHA_7 U1 (C[8], S[7], Y[7], X[7]);
  PureCSA_37_8 U2 (C[38:9], S[37:8], Z[37:8], Y[37:8], X[37:8]);
  UBHA_38 U3 (C[39], S[38], Z[38], Y[38]);
  UB1DCON_39 U4 (S[39], Z[39]);
endmodule

module CSA_39_0_37_4_43_000 (C, S, X, Y, Z);
  output [40:5] C;
  output [43:0] S;
  input [39:0] X;
  input [37:4] Y;
  input [43:7] Z;
  UBCON_3_0 U0 (S[3:0], X[3:0]);
  PureCSHA_6_4 U1 (C[7:5], S[6:4], Y[6:4], X[6:4]);
  PureCSA_37_7 U2 (C[38:8], S[37:7], Z[37:7], Y[37:7], X[37:7]);
  PureCSHA_39_38 U3 (C[40:39], S[39:38], Z[39:38], X[39:38]);
  UBCON_43_40 U4 (S[43:40], Z[43:40]);
endmodule

module CSA_40_7_43_9_43_000 (C, S, X, Y, Z);
  output [44:10] C;
  output [43:7] S;
  input [40:7] X;
  input [43:9] Y;
  input [43:12] Z;
  UBCON_8_7 U0 (S[8:7], X[8:7]);
  PureCSHA_11_9 U1 (C[12:10], S[11:9], Y[11:9], X[11:9]);
  PureCSA_40_12 U2 (C[41:13], S[40:12], Z[40:12], Y[40:12], X[40:12]);
  PureCSHA_43_41 U3 (C[44:42], S[43:41], Z[43:41], Y[43:41]);
endmodule

module CSA_40_9_41_10_42000 (C, S, X, Y, Z);
  output [42:11] C;
  output [42:9] S;
  input [40:9] X;
  input [41:10] Y;
  input [42:11] Z;
  UB1DCON_9 U0 (S[9], X[9]);
  UBHA_10 U1 (C[11], S[10], Y[10], X[10]);
  PureCSA_40_11 U2 (C[41:12], S[40:11], Z[40:11], Y[40:11], X[40:11]);
  UBHA_41 U3 (C[42], S[41], Z[41], Y[41]);
  UB1DCON_42 U4 (S[42], Z[42]);
endmodule

module CSA_42_9_42_11_43000 (C, S, X, Y, Z);
  output [43:12] C;
  output [43:9] S;
  input [42:9] X;
  input [42:11] Y;
  input [43:12] Z;
  UBCON_10_9 U0 (S[10:9], X[10:9]);
  UBHA_11 U1 (C[12], S[11], Y[11], X[11]);
  PureCSA_42_12 U2 (C[43:13], S[42:12], Z[42:12], Y[42:12], X[42:12]);
  UB1DCON_43 U3 (S[43], Z[43]);
endmodule

module CSA_43_0_40_5_49_000 (C, S, X, Y, Z);
  output [44:6] C;
  output [49:0] S;
  input [43:0] X;
  input [40:5] Y;
  input [49:10] Z;
  UBCON_4_0 U0 (S[4:0], X[4:0]);
  PureCSHA_9_5 U1 (C[10:6], S[9:5], Y[9:5], X[9:5]);
  PureCSA_40_10 U2 (C[41:11], S[40:10], Z[40:10], Y[40:10], X[40:10]);
  PureCSHA_43_41 U3 (C[44:42], S[43:41], Z[43:41], X[43:41]);
  UBCON_49_44 U4 (S[49:44], Z[49:44]);
endmodule

module CSA_44_10_49_13_4000 (C, S, X, Y, Z);
  output [48:14] C;
  output [49:10] S;
  input [44:10] X;
  input [49:13] Y;
  input [47:16] Z;
  UBCON_12_10 U0 (S[12:10], X[12:10]);
  PureCSHA_15_13 U1 (C[16:14], S[15:13], Y[15:13], X[15:13]);
  PureCSA_44_16 U2 (C[45:17], S[44:16], Z[44:16], Y[44:16], X[44:16]);
  PureCSHA_47_45 U3 (C[48:46], S[47:45], Y[47:45], Z[47:45]);
  UBCON_49_48 U4 (S[49:48], Y[49:48]);
endmodule

module CSA_44_13_45_14_4000 (C, S, X, Y, Z);
  output [46:15] C;
  output [46:13] S;
  input [44:13] X;
  input [45:14] Y;
  input [46:15] Z;
  UB1DCON_13 U0 (S[13], X[13]);
  UBHA_14 U1 (C[15], S[14], Y[14], X[14]);
  PureCSA_44_15 U2 (C[45:16], S[44:15], Z[44:15], Y[44:15], X[44:15]);
  UBHA_45 U3 (C[46], S[45], Z[45], Y[45]);
  UB1DCON_46 U4 (S[46], Z[46]);
endmodule

module CSA_46_13_46_15_4000 (C, S, X, Y, Z);
  output [47:16] C;
  output [49:13] S;
  input [46:13] X;
  input [46:15] Y;
  input [49:16] Z;
  UBCON_14_13 U0 (S[14:13], X[14:13]);
  UBHA_15 U1 (C[16], S[15], Y[15], X[15]);
  PureCSA_46_16 U2 (C[47:17], S[46:16], Z[46:16], Y[46:16], X[46:16]);
  UBCON_49_47 U3 (S[49:47], Z[49:47]);
endmodule

module CSA_47_16_48_17_4000 (C, S, X, Y, Z);
  output [49:18] C;
  output [49:16] S;
  input [47:16] X;
  input [48:17] Y;
  input [49:18] Z;
  UB1DCON_16 U0 (S[16], X[16]);
  UBHA_17 U1 (C[18], S[17], Y[17], X[17]);
  PureCSA_47_18 U2 (C[48:19], S[47:18], Z[47:18], Y[47:18], X[47:18]);
  UBHA_48 U3 (C[49], S[48], Z[48], Y[48]);
  UB1DCON_49 U4 (S[49], Z[49]);
endmodule

module CSA_48_14_58_18_5000 (C, S, X, Y, Z);
  output [55:19] C;
  output [58:14] S;
  input [48:14] X;
  input [58:18] Y;
  input [54:21] Z;
  UBCON_17_14 U0 (S[17:14], X[17:14]);
  PureCSHA_20_18 U1 (C[21:19], S[20:18], Y[20:18], X[20:18]);
  PureCSA_48_21 U2 (C[49:22], S[48:21], Z[48:21], Y[48:21], X[48:21]);
  PureCSHA_54_49 U3 (C[55:50], S[54:49], Y[54:49], Z[54:49]);
  UBCON_58_55 U4 (S[58:55], Y[58:55]);
endmodule

module CSA_49_0_44_6_58_000 (C, S, X, Y, Z);
  output [50:7] C;
  output [58:0] S;
  input [49:0] X;
  input [44:6] Y;
  input [58:14] Z;
  UBCON_5_0 U0 (S[5:0], X[5:0]);
  PureCSHA_13_6 U1 (C[14:7], S[13:6], Y[13:6], X[13:6]);
  PureCSA_44_14 U2 (C[45:15], S[44:14], Z[44:14], Y[44:14], X[44:14]);
  PureCSHA_49_45 U3 (C[50:46], S[49:45], Z[49:45], X[49:45]);
  UBCON_58_50 U4 (S[58:50], Z[58:50]);
endmodule

module CSA_49_18_52_19_5000 (C, S, X, Y, Z);
  output [53:20] C;
  output [52:18] S;
  input [49:18] X;
  input [52:19] Y;
  input [52:21] Z;
  UB1DCON_18 U0 (S[18], X[18]);
  PureCSHA_20_19 U1 (C[21:20], S[20:19], Y[20:19], X[20:19]);
  PureCSA_49_21 U2 (C[50:22], S[49:21], Z[49:21], Y[49:21], X[49:21]);
  PureCSHA_52_50 U3 (C[53:51], S[52:50], Z[52:50], Y[52:50]);
endmodule

module CSA_50_19_51_20_5000 (C, S, X, Y, Z);
  output [52:21] C;
  output [52:19] S;
  input [50:19] X;
  input [51:20] Y;
  input [52:21] Z;
  UB1DCON_19 U0 (S[19], X[19]);
  UBHA_20 U1 (C[21], S[20], Y[20], X[20]);
  PureCSA_50_21 U2 (C[51:22], S[50:21], Z[50:21], Y[50:21], X[50:21]);
  UBHA_51 U3 (C[52], S[51], Z[51], Y[51]);
  UB1DCON_52 U4 (S[52], Z[52]);
endmodule

module CSA_52_18_53_20_5000 (C, S, X, Y, Z);
  output [54:21] C;
  output [58:18] S;
  input [52:18] X;
  input [53:20] Y;
  input [58:22] Z;
  UBCON_19_18 U0 (S[19:18], X[19:18]);
  PureCSHA_21_20 U1 (C[22:21], S[21:20], Y[21:20], X[21:20]);
  PureCSA_52_22 U2 (C[53:23], S[52:22], Z[52:22], Y[52:22], X[52:22]);
  UBHA_53 U3 (C[54], S[53], Z[53], Y[53]);
  UBCON_58_54 U4 (S[58:54], Z[58:54]);
endmodule

module CSA_53_22_54_23_5000 (C, S, X, Y, Z);
  output [55:24] C;
  output [55:22] S;
  input [53:22] X;
  input [54:23] Y;
  input [55:24] Z;
  UB1DCON_22 U0 (S[22], X[22]);
  UBHA_23 U1 (C[24], S[23], Y[23], X[23]);
  PureCSA_53_24 U2 (C[54:25], S[53:24], Z[53:24], Y[53:24], X[53:24]);
  UBHA_54 U3 (C[55], S[54], Z[54], Y[54]);
  UB1DCON_55 U4 (S[55], Z[55]);
endmodule

module CSA_55_19_62_25_6000 (C, S, X, Y, Z);
  output [63:26] C;
  output [63:19] S;
  input [55:19] X;
  input [62:25] Y;
  input [63:29] Z;
  UBCON_24_19 U0 (S[24:19], X[24:19]);
  PureCSHA_28_25 U1 (C[29:26], S[28:25], Y[28:25], X[28:25]);
  PureCSA_55_29 U2 (C[56:30], S[55:29], Z[55:29], Y[55:29], X[55:29]);
  PureCSHA_62_56 U3 (C[63:57], S[62:56], Z[62:56], Y[62:56]);
  UB1DCON_63 U4 (S[63], Z[63]);
endmodule

module CSA_55_22_55_24_5000 (C, S, X, Y, Z);
  output [56:25] C;
  output [58:22] S;
  input [55:22] X;
  input [55:24] Y;
  input [58:25] Z;
  UBCON_23_22 U0 (S[23:22], X[23:22]);
  UBHA_24 U1 (C[25], S[24], Y[24], X[24]);
  PureCSA_55_25 U2 (C[56:26], S[55:25], Z[55:25], Y[55:25], X[55:25]);
  UBCON_58_56 U3 (S[58:56], Z[58:56]);
endmodule

module CSA_56_25_57_26_5000 (C, S, X, Y, Z);
  output [58:27] C;
  output [58:25] S;
  input [56:25] X;
  input [57:26] Y;
  input [58:27] Z;
  UB1DCON_25 U0 (S[25], X[25]);
  UBHA_26 U1 (C[27], S[26], Y[26], X[26]);
  PureCSA_56_27 U2 (C[57:28], S[56:27], Z[56:27], Y[56:27], X[56:27]);
  UBHA_57 U3 (C[58], S[57], Z[57], Y[57]);
  UB1DCON_58 U4 (S[58], Z[58]);
endmodule

module CSA_56_25_61_27_6000 (C, S, X, Y, Z);
  output [62:28] C;
  output [62:25] S;
  input [56:25] X;
  input [61:27] Y;
  input [62:29] Z;
  UBCON_26_25 U0 (S[26:25], X[26:25]);
  PureCSHA_28_27 U1 (C[29:28], S[28:27], Y[28:27], X[28:27]);
  PureCSA_56_29 U2 (C[57:30], S[56:29], Z[56:29], Y[56:29], X[56:29]);
  PureCSHA_61_57 U3 (C[62:58], S[61:57], Z[61:57], Y[61:57]);
  UB1DCON_62 U4 (S[62], Z[62]);
endmodule

module CSA_58_0_50_7_63_000 (C, S, X, Y, Z);
  output [59:8] C;
  output [63:0] S;
  input [58:0] X;
  input [50:7] Y;
  input [63:19] Z;
  UBCON_6_0 U0 (S[6:0], X[6:0]);
  PureCSHA_18_7 U1 (C[19:8], S[18:7], Y[18:7], X[18:7]);
  PureCSA_50_19 U2 (C[51:20], S[50:19], Z[50:19], Y[50:19], X[50:19]);
  PureCSHA_58_51 U3 (C[59:52], S[58:51], Z[58:51], X[58:51]);
  UBCON_63_59 U4 (S[63:59], Z[63:59]);
endmodule

module CSA_58_27_61_28_6000 (C, S, X, Y, Z);
  output [62:29] C;
  output [61:27] S;
  input [58:27] X;
  input [61:28] Y;
  input [61:30] Z;
  UB1DCON_27 U0 (S[27], X[27]);
  PureCSHA_29_28 U1 (C[30:29], S[29:28], Y[29:28], X[29:28]);
  PureCSA_58_30 U2 (C[59:31], S[58:30], Z[58:30], Y[58:30], X[58:30]);
  PureCSHA_61_59 U3 (C[62:60], S[61:59], Z[61:59], Y[61:59]);
endmodule

module CSA_59_28_60_29_6000 (C, S, X, Y, Z);
  output [61:30] C;
  output [61:28] S;
  input [59:28] X;
  input [60:29] Y;
  input [61:30] Z;
  UB1DCON_28 U0 (S[28], X[28]);
  UBHA_29 U1 (C[30], S[29], Y[29], X[29]);
  PureCSA_59_30 U2 (C[60:31], S[59:30], Z[59:30], Y[59:30], X[59:30]);
  UBHA_60 U3 (C[61], S[60], Z[60], Y[60]);
  UB1DCON_61 U4 (S[61], Z[61]);
endmodule

module CSA_62_25_62_28_6000 (C, S, X, Y, Z);
  output [63:29] C;
  output [62:25] S;
  input [62:25] X;
  input [62:28] Y;
  input [62:31] Z;
  UBCON_27_25 U0 (S[27:25], X[27:25]);
  PureCSHA_30_28 U1 (C[31:29], S[30:28], Y[30:28], X[30:28]);
  PureCSA_62_31 U2 (C[63:32], S[62:31], Z[62:31], Y[62:31], X[62:31]);
endmodule

module CSA_63_0_59_8_63_000 (C, S, X, Y, Z);
  output [64:9] C;
  output [63:0] S;
  input [63:0] X;
  input [59:8] Y;
  input [63:26] Z;
  UBCON_7_0 U0 (S[7:0], X[7:0]);
  PureCSHA_25_8 U1 (C[26:9], S[25:8], Y[25:8], X[25:8]);
  PureCSA_59_26 U2 (C[60:27], S[59:26], Z[59:26], Y[59:26], X[59:26]);
  PureCSHA_63_60 U3 (C[64:61], S[63:60], Z[63:60], X[63:60]);
endmodule

module MultTC_STD_WAL_KS000 (P, IN1, IN2, clk, rst);

  input clk, rst;

  output [66:0] P;
  input [31:0] IN1;
  input [31:0] IN2;
  wire [32:0] PP0;
  wire [32:1] PP1;
  wire [41:10] PP10;
  wire [42:11] PP11;
  wire [43:12] PP12;
  wire [44:13] PP13;
  wire [45:14] PP14;
  wire [46:15] PP15;
  wire [47:16] PP16;
  wire [48:17] PP17;
  wire [49:18] PP18;
  wire [50:19] PP19;
  wire [33:2] PP2;
  wire [51:20] PP20;
  wire [52:21] PP21;
  wire [53:22] PP22;
  wire [54:23] PP23;
  wire [55:24] PP24;
  wire [56:25] PP25;
  wire [57:26] PP26;
  wire [58:27] PP27;
  wire [59:28] PP28;
  wire [60:29] PP29;
  wire [34:3] PP3;
  wire [61:30] PP30;
  wire [62:31] PP31;
  wire [35:4] PP4;
  wire [36:5] PP5;
  wire [37:6] PP6;
  wire [38:7] PP7;
  wire [39:8] PP8;
  wire [40:9] PP9;
  wire [65:0] P_UB;
  wire [64:9] S1;
  wire [63:0] S2;

  reg [64:9] S1_reg;
  reg [63:0] S2_reg;

  TCPPG_31_0_31_0 U0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, IN1, IN2);
  WLCTR_32_0_32_1_3000 U1 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31);

  // amir
  always @(posedge clk)
  begin
    if(rst) begin
      S1_reg <= 0;
      S2_reg <= 0;
    end
    else
    begin
      S1_reg <= S1;
      S2_reg <= S2;
    end
  end
  // rima

  UBKSA_64_9_63_0 U2 (P_UB, S1_reg, S2_reg);
  UBTCCONV63_65_0 U3 (P, P_UB);
endmodule

module NUBUBCON_61_31 (O, I);
  output [61:31] O;
  input [61:31] I;
  NUBUB1CON_31 U0 (O[31], I[31]);
  NUBUB1CON_32 U1 (O[32], I[32]);
  NUBUB1CON_33 U2 (O[33], I[33]);
  NUBUB1CON_34 U3 (O[34], I[34]);
  NUBUB1CON_35 U4 (O[35], I[35]);
  NUBUB1CON_36 U5 (O[36], I[36]);
  NUBUB1CON_37 U6 (O[37], I[37]);
  NUBUB1CON_38 U7 (O[38], I[38]);
  NUBUB1CON_39 U8 (O[39], I[39]);
  NUBUB1CON_40 U9 (O[40], I[40]);
  NUBUB1CON_41 U10 (O[41], I[41]);
  NUBUB1CON_42 U11 (O[42], I[42]);
  NUBUB1CON_43 U12 (O[43], I[43]);
  NUBUB1CON_44 U13 (O[44], I[44]);
  NUBUB1CON_45 U14 (O[45], I[45]);
  NUBUB1CON_46 U15 (O[46], I[46]);
  NUBUB1CON_47 U16 (O[47], I[47]);
  NUBUB1CON_48 U17 (O[48], I[48]);
  NUBUB1CON_49 U18 (O[49], I[49]);
  NUBUB1CON_50 U19 (O[50], I[50]);
  NUBUB1CON_51 U20 (O[51], I[51]);
  NUBUB1CON_52 U21 (O[52], I[52]);
  NUBUB1CON_53 U22 (O[53], I[53]);
  NUBUB1CON_54 U23 (O[54], I[54]);
  NUBUB1CON_55 U24 (O[55], I[55]);
  NUBUB1CON_56 U25 (O[56], I[56]);
  NUBUB1CON_57 U26 (O[57], I[57]);
  NUBUB1CON_58 U27 (O[58], I[58]);
  NUBUB1CON_59 U28 (O[59], I[59]);
  NUBUB1CON_60 U29 (O[60], I[60]);
  NUBUB1CON_61 U30 (O[61], I[61]);
endmodule

module PureCSA_32_2 (C, S, X, Y, Z);
  output [33:3] C;
  output [32:2] S;
  input [32:2] X;
  input [32:2] Y;
  input [32:2] Z;
  UBFA_2 U0 (C[3], S[2], X[2], Y[2], Z[2]);
  UBFA_3 U1 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U2 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U3 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U4 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U5 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U6 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U7 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U8 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U9 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U10 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U11 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U12 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U13 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U14 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U15 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U16 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U17 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U18 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U19 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U20 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U21 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U22 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U23 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U24 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U25 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U26 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U27 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U28 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U29 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U30 (C[33], S[32], X[32], Y[32], Z[32]);
endmodule

module PureCSA_33_3 (C, S, X, Y, Z);
  output [34:4] C;
  output [33:3] S;
  input [33:3] X;
  input [33:3] Y;
  input [33:3] Z;
  UBFA_3 U0 (C[4], S[3], X[3], Y[3], Z[3]);
  UBFA_4 U1 (C[5], S[4], X[4], Y[4], Z[4]);
  UBFA_5 U2 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U3 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U4 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U5 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U6 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U7 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U8 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U9 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U10 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U11 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U12 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U13 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U14 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U15 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U16 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U17 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U18 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U19 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U20 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U21 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U22 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U23 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U24 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U25 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U26 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U27 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U28 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U29 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U30 (C[34], S[33], X[33], Y[33], Z[33]);
endmodule

module PureCSA_34_5 (C, S, X, Y, Z);
  output [35:6] C;
  output [34:5] S;
  input [34:5] X;
  input [34:5] Y;
  input [34:5] Z;
  UBFA_5 U0 (C[6], S[5], X[5], Y[5], Z[5]);
  UBFA_6 U1 (C[7], S[6], X[6], Y[6], Z[6]);
  UBFA_7 U2 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U3 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U4 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U5 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U6 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U7 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U8 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U9 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U10 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U11 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U12 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U13 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U14 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U15 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U16 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U17 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U18 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U19 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U20 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U21 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U22 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U23 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U24 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U25 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U26 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U27 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U28 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U29 (C[35], S[34], X[34], Y[34], Z[34]);
endmodule

module PureCSA_36_8 (C, S, X, Y, Z);
  output [37:9] C;
  output [36:8] S;
  input [36:8] X;
  input [36:8] Y;
  input [36:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U12 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U13 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U14 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U15 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U16 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U17 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U18 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U19 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U20 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U21 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U22 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U23 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U24 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U25 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U26 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U27 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U28 (C[37], S[36], X[36], Y[36], Z[36]);
endmodule

module PureCSA_37_7 (C, S, X, Y, Z);
  output [38:8] C;
  output [37:7] S;
  input [37:7] X;
  input [37:7] Y;
  input [37:7] Z;
  UBFA_7 U0 (C[8], S[7], X[7], Y[7], Z[7]);
  UBFA_8 U1 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U2 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U3 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U4 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U5 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U6 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U7 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U8 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U9 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U10 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U11 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U12 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U13 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U14 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U15 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U16 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U17 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U18 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U19 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U20 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U21 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U22 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U23 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U24 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U25 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U26 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U27 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U28 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U29 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U30 (C[38], S[37], X[37], Y[37], Z[37]);
endmodule

module PureCSA_37_8 (C, S, X, Y, Z);
  output [38:9] C;
  output [37:8] S;
  input [37:8] X;
  input [37:8] Y;
  input [37:8] Z;
  UBFA_8 U0 (C[9], S[8], X[8], Y[8], Z[8]);
  UBFA_9 U1 (C[10], S[9], X[9], Y[9], Z[9]);
  UBFA_10 U2 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U3 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U4 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U5 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U6 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U7 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U8 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U9 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U10 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U11 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U12 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U13 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U14 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U15 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U16 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U17 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U18 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U19 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U20 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U21 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U22 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U23 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U24 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U25 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U26 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U27 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U28 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U29 (C[38], S[37], X[37], Y[37], Z[37]);
endmodule

module PureCSA_40_10 (C, S, X, Y, Z);
  output [41:11] C;
  output [40:10] S;
  input [40:10] X;
  input [40:10] Y;
  input [40:10] Z;
  UBFA_10 U0 (C[11], S[10], X[10], Y[10], Z[10]);
  UBFA_11 U1 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U2 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U3 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U4 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U5 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U6 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U7 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U8 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U9 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U10 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U11 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U12 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U13 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U14 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U15 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U16 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U17 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U18 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U19 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U20 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U21 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U22 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U23 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U24 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U25 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U26 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U27 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U28 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U29 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U30 (C[41], S[40], X[40], Y[40], Z[40]);
endmodule

module PureCSA_40_11 (C, S, X, Y, Z);
  output [41:12] C;
  output [40:11] S;
  input [40:11] X;
  input [40:11] Y;
  input [40:11] Z;
  UBFA_11 U0 (C[12], S[11], X[11], Y[11], Z[11]);
  UBFA_12 U1 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U2 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U3 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U4 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U5 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U6 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U7 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U8 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U9 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U10 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U11 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U12 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U13 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U14 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U15 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U16 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U17 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U18 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U19 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U20 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U21 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U22 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U23 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U24 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U25 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U26 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U27 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U28 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U29 (C[41], S[40], X[40], Y[40], Z[40]);
endmodule

module PureCSA_40_12 (C, S, X, Y, Z);
  output [41:13] C;
  output [40:12] S;
  input [40:12] X;
  input [40:12] Y;
  input [40:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U12 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U13 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U14 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U15 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U16 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U17 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U18 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U19 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U20 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U21 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U22 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U23 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U24 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U25 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U26 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U27 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U28 (C[41], S[40], X[40], Y[40], Z[40]);
endmodule

module PureCSA_42_12 (C, S, X, Y, Z);
  output [43:13] C;
  output [42:12] S;
  input [42:12] X;
  input [42:12] Y;
  input [42:12] Z;
  UBFA_12 U0 (C[13], S[12], X[12], Y[12], Z[12]);
  UBFA_13 U1 (C[14], S[13], X[13], Y[13], Z[13]);
  UBFA_14 U2 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U3 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U4 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U5 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U6 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U7 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U8 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U9 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U10 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U11 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U12 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U13 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U14 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U15 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U16 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U17 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U18 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U19 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U20 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U21 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U22 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U23 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U24 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U25 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U26 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U27 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U28 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U29 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U30 (C[43], S[42], X[42], Y[42], Z[42]);
endmodule

module PureCSA_44_14 (C, S, X, Y, Z);
  output [45:15] C;
  output [44:14] S;
  input [44:14] X;
  input [44:14] Y;
  input [44:14] Z;
  UBFA_14 U0 (C[15], S[14], X[14], Y[14], Z[14]);
  UBFA_15 U1 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U2 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U3 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U4 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U5 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U6 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U7 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U8 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U9 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U10 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U11 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U12 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U13 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U14 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U15 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U16 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U17 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U18 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U19 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U20 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U21 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U22 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U23 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U24 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U25 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U26 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U27 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U28 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U29 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U30 (C[45], S[44], X[44], Y[44], Z[44]);
endmodule

module PureCSA_44_15 (C, S, X, Y, Z);
  output [45:16] C;
  output [44:15] S;
  input [44:15] X;
  input [44:15] Y;
  input [44:15] Z;
  UBFA_15 U0 (C[16], S[15], X[15], Y[15], Z[15]);
  UBFA_16 U1 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U2 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U3 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U4 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U5 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U6 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U7 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U8 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U9 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U10 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U11 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U12 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U13 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U14 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U15 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U16 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U17 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U18 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U19 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U20 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U21 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U22 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U23 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U24 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U25 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U26 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U27 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U28 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U29 (C[45], S[44], X[44], Y[44], Z[44]);
endmodule

module PureCSA_44_16 (C, S, X, Y, Z);
  output [45:17] C;
  output [44:16] S;
  input [44:16] X;
  input [44:16] Y;
  input [44:16] Z;
  UBFA_16 U0 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U1 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U2 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U3 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U4 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U5 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U6 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U7 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U8 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U9 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U10 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U11 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U12 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U13 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U14 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U15 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U16 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U17 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U18 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U19 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U20 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U21 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U22 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U23 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U24 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U25 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U26 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U27 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U28 (C[45], S[44], X[44], Y[44], Z[44]);
endmodule

module PureCSA_46_16 (C, S, X, Y, Z);
  output [47:17] C;
  output [46:16] S;
  input [46:16] X;
  input [46:16] Y;
  input [46:16] Z;
  UBFA_16 U0 (C[17], S[16], X[16], Y[16], Z[16]);
  UBFA_17 U1 (C[18], S[17], X[17], Y[17], Z[17]);
  UBFA_18 U2 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U3 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U4 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U5 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U6 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U7 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U8 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U9 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U10 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U11 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U12 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U13 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U14 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U15 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U16 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U17 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U18 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U19 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U20 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U21 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U22 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U23 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U24 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U25 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U26 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U27 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U28 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U29 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U30 (C[47], S[46], X[46], Y[46], Z[46]);
endmodule

module PureCSA_47_18 (C, S, X, Y, Z);
  output [48:19] C;
  output [47:18] S;
  input [47:18] X;
  input [47:18] Y;
  input [47:18] Z;
  UBFA_18 U0 (C[19], S[18], X[18], Y[18], Z[18]);
  UBFA_19 U1 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U2 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U3 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U4 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U5 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U6 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U7 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U8 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U9 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U10 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U11 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U12 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U13 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U14 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U15 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U16 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U17 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U18 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U19 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U20 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U21 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U22 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U23 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U24 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U25 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U26 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U27 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U28 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U29 (C[48], S[47], X[47], Y[47], Z[47]);
endmodule

module PureCSA_48_21 (C, S, X, Y, Z);
  output [49:22] C;
  output [48:21] S;
  input [48:21] X;
  input [48:21] Y;
  input [48:21] Z;
  UBFA_21 U0 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U1 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U2 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U3 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U4 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U5 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U6 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U7 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U8 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U9 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U10 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U11 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U12 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U13 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U14 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U15 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U16 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U17 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U18 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U19 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U20 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U21 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U22 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U23 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U24 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U25 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U26 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U27 (C[49], S[48], X[48], Y[48], Z[48]);
endmodule

module PureCSA_49_21 (C, S, X, Y, Z);
  output [50:22] C;
  output [49:21] S;
  input [49:21] X;
  input [49:21] Y;
  input [49:21] Z;
  UBFA_21 U0 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U1 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U2 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U3 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U4 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U5 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U6 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U7 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U8 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U9 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U10 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U11 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U12 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U13 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U14 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U15 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U16 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U17 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U18 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U19 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U20 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U21 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U22 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U23 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U24 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U25 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U26 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U27 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U28 (C[50], S[49], X[49], Y[49], Z[49]);
endmodule

module PureCSA_50_19 (C, S, X, Y, Z);
  output [51:20] C;
  output [50:19] S;
  input [50:19] X;
  input [50:19] Y;
  input [50:19] Z;
  UBFA_19 U0 (C[20], S[19], X[19], Y[19], Z[19]);
  UBFA_20 U1 (C[21], S[20], X[20], Y[20], Z[20]);
  UBFA_21 U2 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U3 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U4 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U5 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U6 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U7 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U8 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U9 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U10 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U11 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U12 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U13 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U14 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U15 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U16 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U17 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U18 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U19 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U20 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U21 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U22 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U23 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U24 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U25 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U26 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U27 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U28 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U29 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U30 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U31 (C[51], S[50], X[50], Y[50], Z[50]);
endmodule

module PureCSA_50_21 (C, S, X, Y, Z);
  output [51:22] C;
  output [50:21] S;
  input [50:21] X;
  input [50:21] Y;
  input [50:21] Z;
  UBFA_21 U0 (C[22], S[21], X[21], Y[21], Z[21]);
  UBFA_22 U1 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U2 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U3 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U4 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U5 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U6 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U7 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U8 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U9 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U10 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U11 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U12 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U13 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U14 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U15 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U16 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U17 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U18 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U19 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U20 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U21 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U22 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U23 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U24 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U25 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U26 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U27 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U28 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U29 (C[51], S[50], X[50], Y[50], Z[50]);
endmodule

module PureCSA_52_22 (C, S, X, Y, Z);
  output [53:23] C;
  output [52:22] S;
  input [52:22] X;
  input [52:22] Y;
  input [52:22] Z;
  UBFA_22 U0 (C[23], S[22], X[22], Y[22], Z[22]);
  UBFA_23 U1 (C[24], S[23], X[23], Y[23], Z[23]);
  UBFA_24 U2 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U3 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U4 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U5 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U6 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U7 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U8 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U9 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U10 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U11 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U12 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U13 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U14 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U15 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U16 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U17 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U18 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U19 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U20 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U21 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U22 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U23 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U24 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U25 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U26 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U27 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U28 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U29 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U30 (C[53], S[52], X[52], Y[52], Z[52]);
endmodule

module PureCSA_53_24 (C, S, X, Y, Z);
  output [54:25] C;
  output [53:24] S;
  input [53:24] X;
  input [53:24] Y;
  input [53:24] Z;
  UBFA_24 U0 (C[25], S[24], X[24], Y[24], Z[24]);
  UBFA_25 U1 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U2 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U3 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U4 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U5 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U6 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U7 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U8 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U9 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U10 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U11 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U12 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U13 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U14 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U15 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U16 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U17 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U18 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U19 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U20 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U21 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U22 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U23 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U24 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U25 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U26 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U27 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U28 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U29 (C[54], S[53], X[53], Y[53], Z[53]);
endmodule

module PureCSA_55_25 (C, S, X, Y, Z);
  output [56:26] C;
  output [55:25] S;
  input [55:25] X;
  input [55:25] Y;
  input [55:25] Z;
  UBFA_25 U0 (C[26], S[25], X[25], Y[25], Z[25]);
  UBFA_26 U1 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U2 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U3 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U4 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U5 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U6 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U7 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U8 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U9 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U10 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U11 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U12 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U13 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U14 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U15 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U16 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U17 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U18 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U19 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U20 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U21 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U22 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U23 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U24 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U25 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U26 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U27 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U28 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U29 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U30 (C[56], S[55], X[55], Y[55], Z[55]);
endmodule

module PureCSA_55_29 (C, S, X, Y, Z);
  output [56:30] C;
  output [55:29] S;
  input [55:29] X;
  input [55:29] Y;
  input [55:29] Z;
  UBFA_29 U0 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U1 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U2 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U3 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U4 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U5 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U6 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U7 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U8 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U9 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U10 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U11 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U12 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U13 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U14 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U15 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U16 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U17 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U18 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U19 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U20 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U21 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U22 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U23 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U24 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U25 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U26 (C[56], S[55], X[55], Y[55], Z[55]);
endmodule

module PureCSA_56_27 (C, S, X, Y, Z);
  output [57:28] C;
  output [56:27] S;
  input [56:27] X;
  input [56:27] Y;
  input [56:27] Z;
  UBFA_27 U0 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U1 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U2 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U3 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U4 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U5 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U6 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U7 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U8 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U9 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U10 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U11 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U12 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U13 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U14 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U15 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U16 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U17 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U18 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U19 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U20 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U21 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U22 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U23 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U24 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U25 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U26 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U27 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U28 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U29 (C[57], S[56], X[56], Y[56], Z[56]);
endmodule

module PureCSA_56_29 (C, S, X, Y, Z);
  output [57:30] C;
  output [56:29] S;
  input [56:29] X;
  input [56:29] Y;
  input [56:29] Z;
  UBFA_29 U0 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U1 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U2 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U3 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U4 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U5 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U6 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U7 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U8 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U9 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U10 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U11 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U12 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U13 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U14 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U15 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U16 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U17 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U18 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U19 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U20 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U21 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U22 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U23 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U24 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U25 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U26 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U27 (C[57], S[56], X[56], Y[56], Z[56]);
endmodule

module PureCSA_58_30 (C, S, X, Y, Z);
  output [59:31] C;
  output [58:30] S;
  input [58:30] X;
  input [58:30] Y;
  input [58:30] Z;
  UBFA_30 U0 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U1 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U2 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U3 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U4 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U5 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U6 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U7 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U8 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U9 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U10 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U11 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U12 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U13 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U14 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U15 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U16 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U17 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U18 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U19 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U20 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U21 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U22 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U23 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U24 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U25 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U26 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U27 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U28 (C[59], S[58], X[58], Y[58], Z[58]);
endmodule

module PureCSA_59_26 (C, S, X, Y, Z);
  output [60:27] C;
  output [59:26] S;
  input [59:26] X;
  input [59:26] Y;
  input [59:26] Z;
  UBFA_26 U0 (C[27], S[26], X[26], Y[26], Z[26]);
  UBFA_27 U1 (C[28], S[27], X[27], Y[27], Z[27]);
  UBFA_28 U2 (C[29], S[28], X[28], Y[28], Z[28]);
  UBFA_29 U3 (C[30], S[29], X[29], Y[29], Z[29]);
  UBFA_30 U4 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U5 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U6 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U7 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U8 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U9 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U10 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U11 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U12 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U13 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U14 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U15 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U16 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U17 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U18 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U19 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U20 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U21 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U22 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U23 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U24 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U25 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U26 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U27 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U28 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U29 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U30 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U31 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U32 (C[59], S[58], X[58], Y[58], Z[58]);
  UBFA_59 U33 (C[60], S[59], X[59], Y[59], Z[59]);
endmodule

module PureCSA_59_30 (C, S, X, Y, Z);
  output [60:31] C;
  output [59:30] S;
  input [59:30] X;
  input [59:30] Y;
  input [59:30] Z;
  UBFA_30 U0 (C[31], S[30], X[30], Y[30], Z[30]);
  UBFA_31 U1 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U2 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U3 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U4 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U5 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U6 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U7 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U8 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U9 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U10 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U11 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U12 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U13 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U14 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U15 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U16 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U17 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U18 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U19 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U20 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U21 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U22 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U23 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U24 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U25 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U26 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U27 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U28 (C[59], S[58], X[58], Y[58], Z[58]);
  UBFA_59 U29 (C[60], S[59], X[59], Y[59], Z[59]);
endmodule

module PureCSA_62_31 (C, S, X, Y, Z);
  output [63:32] C;
  output [62:31] S;
  input [62:31] X;
  input [62:31] Y;
  input [62:31] Z;
  UBFA_31 U0 (C[32], S[31], X[31], Y[31], Z[31]);
  UBFA_32 U1 (C[33], S[32], X[32], Y[32], Z[32]);
  UBFA_33 U2 (C[34], S[33], X[33], Y[33], Z[33]);
  UBFA_34 U3 (C[35], S[34], X[34], Y[34], Z[34]);
  UBFA_35 U4 (C[36], S[35], X[35], Y[35], Z[35]);
  UBFA_36 U5 (C[37], S[36], X[36], Y[36], Z[36]);
  UBFA_37 U6 (C[38], S[37], X[37], Y[37], Z[37]);
  UBFA_38 U7 (C[39], S[38], X[38], Y[38], Z[38]);
  UBFA_39 U8 (C[40], S[39], X[39], Y[39], Z[39]);
  UBFA_40 U9 (C[41], S[40], X[40], Y[40], Z[40]);
  UBFA_41 U10 (C[42], S[41], X[41], Y[41], Z[41]);
  UBFA_42 U11 (C[43], S[42], X[42], Y[42], Z[42]);
  UBFA_43 U12 (C[44], S[43], X[43], Y[43], Z[43]);
  UBFA_44 U13 (C[45], S[44], X[44], Y[44], Z[44]);
  UBFA_45 U14 (C[46], S[45], X[45], Y[45], Z[45]);
  UBFA_46 U15 (C[47], S[46], X[46], Y[46], Z[46]);
  UBFA_47 U16 (C[48], S[47], X[47], Y[47], Z[47]);
  UBFA_48 U17 (C[49], S[48], X[48], Y[48], Z[48]);
  UBFA_49 U18 (C[50], S[49], X[49], Y[49], Z[49]);
  UBFA_50 U19 (C[51], S[50], X[50], Y[50], Z[50]);
  UBFA_51 U20 (C[52], S[51], X[51], Y[51], Z[51]);
  UBFA_52 U21 (C[53], S[52], X[52], Y[52], Z[52]);
  UBFA_53 U22 (C[54], S[53], X[53], Y[53], Z[53]);
  UBFA_54 U23 (C[55], S[54], X[54], Y[54], Z[54]);
  UBFA_55 U24 (C[56], S[55], X[55], Y[55], Z[55]);
  UBFA_56 U25 (C[57], S[56], X[56], Y[56], Z[56]);
  UBFA_57 U26 (C[58], S[57], X[57], Y[57], Z[57]);
  UBFA_58 U27 (C[59], S[58], X[58], Y[58], Z[58]);
  UBFA_59 U28 (C[60], S[59], X[59], Y[59], Z[59]);
  UBFA_60 U29 (C[61], S[60], X[60], Y[60], Z[60]);
  UBFA_61 U30 (C[62], S[61], X[61], Y[61], Z[61]);
  UBFA_62 U31 (C[63], S[62], X[62], Y[62], Z[62]);
endmodule

module PureCSHA_11_9 (C, S, X, Y);
  output [12:10] C;
  output [11:9] S;
  input [11:9] X;
  input [11:9] Y;
  UBHA_9 U0 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U1 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U2 (C[12], S[11], X[11], Y[11]);
endmodule

module PureCSHA_13_6 (C, S, X, Y);
  output [14:7] C;
  output [13:6] S;
  input [13:6] X;
  input [13:6] Y;
  UBHA_6 U0 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U1 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U2 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U3 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U4 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U5 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U6 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U7 (C[14], S[13], X[13], Y[13]);
endmodule

module PureCSHA_15_13 (C, S, X, Y);
  output [16:14] C;
  output [15:13] S;
  input [15:13] X;
  input [15:13] Y;
  UBHA_13 U0 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U1 (C[15], S[14], X[14], Y[14]);
  UBHA_15 U2 (C[16], S[15], X[15], Y[15]);
endmodule

module PureCSHA_18_7 (C, S, X, Y);
  output [19:8] C;
  output [18:7] S;
  input [18:7] X;
  input [18:7] Y;
  UBHA_7 U0 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U1 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U2 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U3 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U4 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U5 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U6 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U7 (C[15], S[14], X[14], Y[14]);
  UBHA_15 U8 (C[16], S[15], X[15], Y[15]);
  UBHA_16 U9 (C[17], S[16], X[16], Y[16]);
  UBHA_17 U10 (C[18], S[17], X[17], Y[17]);
  UBHA_18 U11 (C[19], S[18], X[18], Y[18]);
endmodule

module PureCSHA_20_18 (C, S, X, Y);
  output [21:19] C;
  output [20:18] S;
  input [20:18] X;
  input [20:18] Y;
  UBHA_18 U0 (C[19], S[18], X[18], Y[18]);
  UBHA_19 U1 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U2 (C[21], S[20], X[20], Y[20]);
endmodule

module PureCSHA_20_19 (C, S, X, Y);
  output [21:20] C;
  output [20:19] S;
  input [20:19] X;
  input [20:19] Y;
  UBHA_19 U0 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U1 (C[21], S[20], X[20], Y[20]);
endmodule

module PureCSHA_21_20 (C, S, X, Y);
  output [22:21] C;
  output [21:20] S;
  input [21:20] X;
  input [21:20] Y;
  UBHA_20 U0 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U1 (C[22], S[21], X[21], Y[21]);
endmodule

module PureCSHA_25_8 (C, S, X, Y);
  output [26:9] C;
  output [25:8] S;
  input [25:8] X;
  input [25:8] Y;
  UBHA_8 U0 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U1 (C[10], S[9], X[9], Y[9]);
  UBHA_10 U2 (C[11], S[10], X[10], Y[10]);
  UBHA_11 U3 (C[12], S[11], X[11], Y[11]);
  UBHA_12 U4 (C[13], S[12], X[12], Y[12]);
  UBHA_13 U5 (C[14], S[13], X[13], Y[13]);
  UBHA_14 U6 (C[15], S[14], X[14], Y[14]);
  UBHA_15 U7 (C[16], S[15], X[15], Y[15]);
  UBHA_16 U8 (C[17], S[16], X[16], Y[16]);
  UBHA_17 U9 (C[18], S[17], X[17], Y[17]);
  UBHA_18 U10 (C[19], S[18], X[18], Y[18]);
  UBHA_19 U11 (C[20], S[19], X[19], Y[19]);
  UBHA_20 U12 (C[21], S[20], X[20], Y[20]);
  UBHA_21 U13 (C[22], S[21], X[21], Y[21]);
  UBHA_22 U14 (C[23], S[22], X[22], Y[22]);
  UBHA_23 U15 (C[24], S[23], X[23], Y[23]);
  UBHA_24 U16 (C[25], S[24], X[24], Y[24]);
  UBHA_25 U17 (C[26], S[25], X[25], Y[25]);
endmodule

module PureCSHA_28_25 (C, S, X, Y);
  output [29:26] C;
  output [28:25] S;
  input [28:25] X;
  input [28:25] Y;
  UBHA_25 U0 (C[26], S[25], X[25], Y[25]);
  UBHA_26 U1 (C[27], S[26], X[26], Y[26]);
  UBHA_27 U2 (C[28], S[27], X[27], Y[27]);
  UBHA_28 U3 (C[29], S[28], X[28], Y[28]);
endmodule

module PureCSHA_28_27 (C, S, X, Y);
  output [29:28] C;
  output [28:27] S;
  input [28:27] X;
  input [28:27] Y;
  UBHA_27 U0 (C[28], S[27], X[27], Y[27]);
  UBHA_28 U1 (C[29], S[28], X[28], Y[28]);
endmodule

module PureCSHA_29_28 (C, S, X, Y);
  output [30:29] C;
  output [29:28] S;
  input [29:28] X;
  input [29:28] Y;
  UBHA_28 U0 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U1 (C[30], S[29], X[29], Y[29]);
endmodule

module PureCSHA_30_28 (C, S, X, Y);
  output [31:29] C;
  output [30:28] S;
  input [30:28] X;
  input [30:28] Y;
  UBHA_28 U0 (C[29], S[28], X[28], Y[28]);
  UBHA_29 U1 (C[30], S[29], X[29], Y[29]);
  UBHA_30 U2 (C[31], S[30], X[30], Y[30]);
endmodule

module PureCSHA_36_35 (C, S, X, Y);
  output [37:36] C;
  output [36:35] S;
  input [36:35] X;
  input [36:35] Y;
  UBHA_35 U0 (C[36], S[35], X[35], Y[35]);
  UBHA_36 U1 (C[37], S[36], X[36], Y[36]);
endmodule

module PureCSHA_39_37 (C, S, X, Y);
  output [40:38] C;
  output [39:37] S;
  input [39:37] X;
  input [39:37] Y;
  UBHA_37 U0 (C[38], S[37], X[37], Y[37]);
  UBHA_38 U1 (C[39], S[38], X[38], Y[38]);
  UBHA_39 U2 (C[40], S[39], X[39], Y[39]);
endmodule

module PureCSHA_39_38 (C, S, X, Y);
  output [40:39] C;
  output [39:38] S;
  input [39:38] X;
  input [39:38] Y;
  UBHA_38 U0 (C[39], S[38], X[38], Y[38]);
  UBHA_39 U1 (C[40], S[39], X[39], Y[39]);
endmodule

module PureCSHA_43_41 (C, S, X, Y);
  output [44:42] C;
  output [43:41] S;
  input [43:41] X;
  input [43:41] Y;
  UBHA_41 U0 (C[42], S[41], X[41], Y[41]);
  UBHA_42 U1 (C[43], S[42], X[42], Y[42]);
  UBHA_43 U2 (C[44], S[43], X[43], Y[43]);
endmodule

module PureCSHA_47_45 (C, S, X, Y);
  output [48:46] C;
  output [47:45] S;
  input [47:45] X;
  input [47:45] Y;
  UBHA_45 U0 (C[46], S[45], X[45], Y[45]);
  UBHA_46 U1 (C[47], S[46], X[46], Y[46]);
  UBHA_47 U2 (C[48], S[47], X[47], Y[47]);
endmodule

module PureCSHA_49_45 (C, S, X, Y);
  output [50:46] C;
  output [49:45] S;
  input [49:45] X;
  input [49:45] Y;
  UBHA_45 U0 (C[46], S[45], X[45], Y[45]);
  UBHA_46 U1 (C[47], S[46], X[46], Y[46]);
  UBHA_47 U2 (C[48], S[47], X[47], Y[47]);
  UBHA_48 U3 (C[49], S[48], X[48], Y[48]);
  UBHA_49 U4 (C[50], S[49], X[49], Y[49]);
endmodule

module PureCSHA_4_3 (C, S, X, Y);
  output [5:4] C;
  output [4:3] S;
  input [4:3] X;
  input [4:3] Y;
  UBHA_3 U0 (C[4], S[3], X[3], Y[3]);
  UBHA_4 U1 (C[5], S[4], X[4], Y[4]);
endmodule

module PureCSHA_52_50 (C, S, X, Y);
  output [53:51] C;
  output [52:50] S;
  input [52:50] X;
  input [52:50] Y;
  UBHA_50 U0 (C[51], S[50], X[50], Y[50]);
  UBHA_51 U1 (C[52], S[51], X[51], Y[51]);
  UBHA_52 U2 (C[53], S[52], X[52], Y[52]);
endmodule

module PureCSHA_54_49 (C, S, X, Y);
  output [55:50] C;
  output [54:49] S;
  input [54:49] X;
  input [54:49] Y;
  UBHA_49 U0 (C[50], S[49], X[49], Y[49]);
  UBHA_50 U1 (C[51], S[50], X[50], Y[50]);
  UBHA_51 U2 (C[52], S[51], X[51], Y[51]);
  UBHA_52 U3 (C[53], S[52], X[52], Y[52]);
  UBHA_53 U4 (C[54], S[53], X[53], Y[53]);
  UBHA_54 U5 (C[55], S[54], X[54], Y[54]);
endmodule

module PureCSHA_58_51 (C, S, X, Y);
  output [59:52] C;
  output [58:51] S;
  input [58:51] X;
  input [58:51] Y;
  UBHA_51 U0 (C[52], S[51], X[51], Y[51]);
  UBHA_52 U1 (C[53], S[52], X[52], Y[52]);
  UBHA_53 U2 (C[54], S[53], X[53], Y[53]);
  UBHA_54 U3 (C[55], S[54], X[54], Y[54]);
  UBHA_55 U4 (C[56], S[55], X[55], Y[55]);
  UBHA_56 U5 (C[57], S[56], X[56], Y[56]);
  UBHA_57 U6 (C[58], S[57], X[57], Y[57]);
  UBHA_58 U7 (C[59], S[58], X[58], Y[58]);
endmodule

module PureCSHA_61_57 (C, S, X, Y);
  output [62:58] C;
  output [61:57] S;
  input [61:57] X;
  input [61:57] Y;
  UBHA_57 U0 (C[58], S[57], X[57], Y[57]);
  UBHA_58 U1 (C[59], S[58], X[58], Y[58]);
  UBHA_59 U2 (C[60], S[59], X[59], Y[59]);
  UBHA_60 U3 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U4 (C[62], S[61], X[61], Y[61]);
endmodule

module PureCSHA_61_59 (C, S, X, Y);
  output [62:60] C;
  output [61:59] S;
  input [61:59] X;
  input [61:59] Y;
  UBHA_59 U0 (C[60], S[59], X[59], Y[59]);
  UBHA_60 U1 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U2 (C[62], S[61], X[61], Y[61]);
endmodule

module PureCSHA_62_56 (C, S, X, Y);
  output [63:57] C;
  output [62:56] S;
  input [62:56] X;
  input [62:56] Y;
  UBHA_56 U0 (C[57], S[56], X[56], Y[56]);
  UBHA_57 U1 (C[58], S[57], X[57], Y[57]);
  UBHA_58 U2 (C[59], S[58], X[58], Y[58]);
  UBHA_59 U3 (C[60], S[59], X[59], Y[59]);
  UBHA_60 U4 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U5 (C[62], S[61], X[61], Y[61]);
  UBHA_62 U6 (C[63], S[62], X[62], Y[62]);
endmodule

module PureCSHA_63_60 (C, S, X, Y);
  output [64:61] C;
  output [63:60] S;
  input [63:60] X;
  input [63:60] Y;
  UBHA_60 U0 (C[61], S[60], X[60], Y[60]);
  UBHA_61 U1 (C[62], S[61], X[61], Y[61]);
  UBHA_62 U2 (C[63], S[62], X[62], Y[62]);
  UBHA_63 U3 (C[64], S[63], X[63], Y[63]);
endmodule

module PureCSHA_6_4 (C, S, X, Y);
  output [7:5] C;
  output [6:4] S;
  input [6:4] X;
  input [6:4] Y;
  UBHA_4 U0 (C[5], S[4], X[4], Y[4]);
  UBHA_5 U1 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U2 (C[7], S[6], X[6], Y[6]);
endmodule

module PureCSHA_7_6 (C, S, X, Y);
  output [8:7] C;
  output [7:6] S;
  input [7:6] X;
  input [7:6] Y;
  UBHA_6 U0 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U1 (C[8], S[7], X[7], Y[7]);
endmodule

module PureCSHA_9_5 (C, S, X, Y);
  output [10:6] C;
  output [9:5] S;
  input [9:5] X;
  input [9:5] Y;
  UBHA_5 U0 (C[6], S[5], X[5], Y[5]);
  UBHA_6 U1 (C[7], S[6], X[6], Y[6]);
  UBHA_7 U2 (C[8], S[7], X[7], Y[7]);
  UBHA_8 U3 (C[9], S[8], X[8], Y[8]);
  UBHA_9 U4 (C[10], S[9], X[9], Y[9]);
endmodule

module TCNVPPG_31_0_31 (O, IN1, IN2);
  output [62:31] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire [61:31] NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UN1BPPG_0_31 U1 (NEG[31], IN1P[0], IN2);
  UN1BPPG_1_31 U2 (NEG[32], IN1P[1], IN2);
  UN1BPPG_2_31 U3 (NEG[33], IN1P[2], IN2);
  UN1BPPG_3_31 U4 (NEG[34], IN1P[3], IN2);
  UN1BPPG_4_31 U5 (NEG[35], IN1P[4], IN2);
  UN1BPPG_5_31 U6 (NEG[36], IN1P[5], IN2);
  UN1BPPG_6_31 U7 (NEG[37], IN1P[6], IN2);
  UN1BPPG_7_31 U8 (NEG[38], IN1P[7], IN2);
  UN1BPPG_8_31 U9 (NEG[39], IN1P[8], IN2);
  UN1BPPG_9_31 U10 (NEG[40], IN1P[9], IN2);
  UN1BPPG_10_31 U11 (NEG[41], IN1P[10], IN2);
  UN1BPPG_11_31 U12 (NEG[42], IN1P[11], IN2);
  UN1BPPG_12_31 U13 (NEG[43], IN1P[12], IN2);
  UN1BPPG_13_31 U14 (NEG[44], IN1P[13], IN2);
  UN1BPPG_14_31 U15 (NEG[45], IN1P[14], IN2);
  UN1BPPG_15_31 U16 (NEG[46], IN1P[15], IN2);
  UN1BPPG_16_31 U17 (NEG[47], IN1P[16], IN2);
  UN1BPPG_17_31 U18 (NEG[48], IN1P[17], IN2);
  UN1BPPG_18_31 U19 (NEG[49], IN1P[18], IN2);
  UN1BPPG_19_31 U20 (NEG[50], IN1P[19], IN2);
  UN1BPPG_20_31 U21 (NEG[51], IN1P[20], IN2);
  UN1BPPG_21_31 U22 (NEG[52], IN1P[21], IN2);
  UN1BPPG_22_31 U23 (NEG[53], IN1P[22], IN2);
  UN1BPPG_23_31 U24 (NEG[54], IN1P[23], IN2);
  UN1BPPG_24_31 U25 (NEG[55], IN1P[24], IN2);
  UN1BPPG_25_31 U26 (NEG[56], IN1P[25], IN2);
  UN1BPPG_26_31 U27 (NEG[57], IN1P[26], IN2);
  UN1BPPG_27_31 U28 (NEG[58], IN1P[27], IN2);
  UN1BPPG_28_31 U29 (NEG[59], IN1P[28], IN2);
  UN1BPPG_29_31 U30 (NEG[60], IN1P[29], IN2);
  UN1BPPG_30_31 U31 (NEG[61], IN1P[30], IN2);
  NUB1BPPG_31_31 U32 (O[62], IN1N, IN2);
  NUBUBCON_61_31 U33 (O[61:31], NEG);
endmodule

module TCPPG_31_0_31_0 (PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31, IN1, IN2);
  output [32:0] PP0;
  output [32:1] PP1;
  output [41:10] PP10;
  output [42:11] PP11;
  output [43:12] PP12;
  output [44:13] PP13;
  output [45:14] PP14;
  output [46:15] PP15;
  output [47:16] PP16;
  output [48:17] PP17;
  output [49:18] PP18;
  output [50:19] PP19;
  output [33:2] PP2;
  output [51:20] PP20;
  output [52:21] PP21;
  output [53:22] PP22;
  output [54:23] PP23;
  output [55:24] PP24;
  output [56:25] PP25;
  output [57:26] PP26;
  output [58:27] PP27;
  output [59:28] PP28;
  output [60:29] PP29;
  output [34:3] PP3;
  output [61:30] PP30;
  output [62:31] PP31;
  output [35:4] PP4;
  output [36:5] PP5;
  output [37:6] PP6;
  output [38:7] PP7;
  output [39:8] PP8;
  output [40:9] PP9;
  input [31:0] IN1;
  input [31:0] IN2;
  wire BIAS;
  wire [30:0] IN2R;
  wire IN2T;
  wire [31:0] W;
  TCDECON_31_0 U0 (IN2T, IN2R, IN2);
  TCUVPPG_31_0_0 U1 (W, IN1, IN2R[0]);
  TCUVPPG_31_0_1 U2 (PP1, IN1, IN2R[1]);
  TCUVPPG_31_0_2 U3 (PP2, IN1, IN2R[2]);
  TCUVPPG_31_0_3 U4 (PP3, IN1, IN2R[3]);
  TCUVPPG_31_0_4 U5 (PP4, IN1, IN2R[4]);
  TCUVPPG_31_0_5 U6 (PP5, IN1, IN2R[5]);
  TCUVPPG_31_0_6 U7 (PP6, IN1, IN2R[6]);
  TCUVPPG_31_0_7 U8 (PP7, IN1, IN2R[7]);
  TCUVPPG_31_0_8 U9 (PP8, IN1, IN2R[8]);
  TCUVPPG_31_0_9 U10 (PP9, IN1, IN2R[9]);
  TCUVPPG_31_0_10 U11 (PP10, IN1, IN2R[10]);
  TCUVPPG_31_0_11 U12 (PP11, IN1, IN2R[11]);
  TCUVPPG_31_0_12 U13 (PP12, IN1, IN2R[12]);
  TCUVPPG_31_0_13 U14 (PP13, IN1, IN2R[13]);
  TCUVPPG_31_0_14 U15 (PP14, IN1, IN2R[14]);
  TCUVPPG_31_0_15 U16 (PP15, IN1, IN2R[15]);
  TCUVPPG_31_0_16 U17 (PP16, IN1, IN2R[16]);
  TCUVPPG_31_0_17 U18 (PP17, IN1, IN2R[17]);
  TCUVPPG_31_0_18 U19 (PP18, IN1, IN2R[18]);
  TCUVPPG_31_0_19 U20 (PP19, IN1, IN2R[19]);
  TCUVPPG_31_0_20 U21 (PP20, IN1, IN2R[20]);
  TCUVPPG_31_0_21 U22 (PP21, IN1, IN2R[21]);
  TCUVPPG_31_0_22 U23 (PP22, IN1, IN2R[22]);
  TCUVPPG_31_0_23 U24 (PP23, IN1, IN2R[23]);
  TCUVPPG_31_0_24 U25 (PP24, IN1, IN2R[24]);
  TCUVPPG_31_0_25 U26 (PP25, IN1, IN2R[25]);
  TCUVPPG_31_0_26 U27 (PP26, IN1, IN2R[26]);
  TCUVPPG_31_0_27 U28 (PP27, IN1, IN2R[27]);
  TCUVPPG_31_0_28 U29 (PP28, IN1, IN2R[28]);
  TCUVPPG_31_0_29 U30 (PP29, IN1, IN2R[29]);
  TCUVPPG_31_0_30 U31 (PP30, IN1, IN2R[30]);
  TCNVPPG_31_0_31 U32 (PP31, IN1, IN2T);
  UBOne_32 U33 (BIAS);
  UBCMBIN_32_32_31_000 U34 (PP0, BIAS, W);
endmodule

module TCUVPPG_31_0_0 (O, IN1, IN2);
  output [31:0] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_0 U1 (O[0], IN1P[0], IN2);
  UB1BPPG_1_0 U2 (O[1], IN1P[1], IN2);
  UB1BPPG_2_0 U3 (O[2], IN1P[2], IN2);
  UB1BPPG_3_0 U4 (O[3], IN1P[3], IN2);
  UB1BPPG_4_0 U5 (O[4], IN1P[4], IN2);
  UB1BPPG_5_0 U6 (O[5], IN1P[5], IN2);
  UB1BPPG_6_0 U7 (O[6], IN1P[6], IN2);
  UB1BPPG_7_0 U8 (O[7], IN1P[7], IN2);
  UB1BPPG_8_0 U9 (O[8], IN1P[8], IN2);
  UB1BPPG_9_0 U10 (O[9], IN1P[9], IN2);
  UB1BPPG_10_0 U11 (O[10], IN1P[10], IN2);
  UB1BPPG_11_0 U12 (O[11], IN1P[11], IN2);
  UB1BPPG_12_0 U13 (O[12], IN1P[12], IN2);
  UB1BPPG_13_0 U14 (O[13], IN1P[13], IN2);
  UB1BPPG_14_0 U15 (O[14], IN1P[14], IN2);
  UB1BPPG_15_0 U16 (O[15], IN1P[15], IN2);
  UB1BPPG_16_0 U17 (O[16], IN1P[16], IN2);
  UB1BPPG_17_0 U18 (O[17], IN1P[17], IN2);
  UB1BPPG_18_0 U19 (O[18], IN1P[18], IN2);
  UB1BPPG_19_0 U20 (O[19], IN1P[19], IN2);
  UB1BPPG_20_0 U21 (O[20], IN1P[20], IN2);
  UB1BPPG_21_0 U22 (O[21], IN1P[21], IN2);
  UB1BPPG_22_0 U23 (O[22], IN1P[22], IN2);
  UB1BPPG_23_0 U24 (O[23], IN1P[23], IN2);
  UB1BPPG_24_0 U25 (O[24], IN1P[24], IN2);
  UB1BPPG_25_0 U26 (O[25], IN1P[25], IN2);
  UB1BPPG_26_0 U27 (O[26], IN1P[26], IN2);
  UB1BPPG_27_0 U28 (O[27], IN1P[27], IN2);
  UB1BPPG_28_0 U29 (O[28], IN1P[28], IN2);
  UB1BPPG_29_0 U30 (O[29], IN1P[29], IN2);
  UB1BPPG_30_0 U31 (O[30], IN1P[30], IN2);
  NU1BPPG_31_0 U32 (NEG, IN1N, IN2);
  NUBUB1CON_31 U33 (O[31], NEG);
endmodule

module TCUVPPG_31_0_1 (O, IN1, IN2);
  output [32:1] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_1 U1 (O[1], IN1P[0], IN2);
  UB1BPPG_1_1 U2 (O[2], IN1P[1], IN2);
  UB1BPPG_2_1 U3 (O[3], IN1P[2], IN2);
  UB1BPPG_3_1 U4 (O[4], IN1P[3], IN2);
  UB1BPPG_4_1 U5 (O[5], IN1P[4], IN2);
  UB1BPPG_5_1 U6 (O[6], IN1P[5], IN2);
  UB1BPPG_6_1 U7 (O[7], IN1P[6], IN2);
  UB1BPPG_7_1 U8 (O[8], IN1P[7], IN2);
  UB1BPPG_8_1 U9 (O[9], IN1P[8], IN2);
  UB1BPPG_9_1 U10 (O[10], IN1P[9], IN2);
  UB1BPPG_10_1 U11 (O[11], IN1P[10], IN2);
  UB1BPPG_11_1 U12 (O[12], IN1P[11], IN2);
  UB1BPPG_12_1 U13 (O[13], IN1P[12], IN2);
  UB1BPPG_13_1 U14 (O[14], IN1P[13], IN2);
  UB1BPPG_14_1 U15 (O[15], IN1P[14], IN2);
  UB1BPPG_15_1 U16 (O[16], IN1P[15], IN2);
  UB1BPPG_16_1 U17 (O[17], IN1P[16], IN2);
  UB1BPPG_17_1 U18 (O[18], IN1P[17], IN2);
  UB1BPPG_18_1 U19 (O[19], IN1P[18], IN2);
  UB1BPPG_19_1 U20 (O[20], IN1P[19], IN2);
  UB1BPPG_20_1 U21 (O[21], IN1P[20], IN2);
  UB1BPPG_21_1 U22 (O[22], IN1P[21], IN2);
  UB1BPPG_22_1 U23 (O[23], IN1P[22], IN2);
  UB1BPPG_23_1 U24 (O[24], IN1P[23], IN2);
  UB1BPPG_24_1 U25 (O[25], IN1P[24], IN2);
  UB1BPPG_25_1 U26 (O[26], IN1P[25], IN2);
  UB1BPPG_26_1 U27 (O[27], IN1P[26], IN2);
  UB1BPPG_27_1 U28 (O[28], IN1P[27], IN2);
  UB1BPPG_28_1 U29 (O[29], IN1P[28], IN2);
  UB1BPPG_29_1 U30 (O[30], IN1P[29], IN2);
  UB1BPPG_30_1 U31 (O[31], IN1P[30], IN2);
  NU1BPPG_31_1 U32 (NEG, IN1N, IN2);
  NUBUB1CON_32 U33 (O[32], NEG);
endmodule

module TCUVPPG_31_0_10 (O, IN1, IN2);
  output [41:10] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_10 U1 (O[10], IN1P[0], IN2);
  UB1BPPG_1_10 U2 (O[11], IN1P[1], IN2);
  UB1BPPG_2_10 U3 (O[12], IN1P[2], IN2);
  UB1BPPG_3_10 U4 (O[13], IN1P[3], IN2);
  UB1BPPG_4_10 U5 (O[14], IN1P[4], IN2);
  UB1BPPG_5_10 U6 (O[15], IN1P[5], IN2);
  UB1BPPG_6_10 U7 (O[16], IN1P[6], IN2);
  UB1BPPG_7_10 U8 (O[17], IN1P[7], IN2);
  UB1BPPG_8_10 U9 (O[18], IN1P[8], IN2);
  UB1BPPG_9_10 U10 (O[19], IN1P[9], IN2);
  UB1BPPG_10_10 U11 (O[20], IN1P[10], IN2);
  UB1BPPG_11_10 U12 (O[21], IN1P[11], IN2);
  UB1BPPG_12_10 U13 (O[22], IN1P[12], IN2);
  UB1BPPG_13_10 U14 (O[23], IN1P[13], IN2);
  UB1BPPG_14_10 U15 (O[24], IN1P[14], IN2);
  UB1BPPG_15_10 U16 (O[25], IN1P[15], IN2);
  UB1BPPG_16_10 U17 (O[26], IN1P[16], IN2);
  UB1BPPG_17_10 U18 (O[27], IN1P[17], IN2);
  UB1BPPG_18_10 U19 (O[28], IN1P[18], IN2);
  UB1BPPG_19_10 U20 (O[29], IN1P[19], IN2);
  UB1BPPG_20_10 U21 (O[30], IN1P[20], IN2);
  UB1BPPG_21_10 U22 (O[31], IN1P[21], IN2);
  UB1BPPG_22_10 U23 (O[32], IN1P[22], IN2);
  UB1BPPG_23_10 U24 (O[33], IN1P[23], IN2);
  UB1BPPG_24_10 U25 (O[34], IN1P[24], IN2);
  UB1BPPG_25_10 U26 (O[35], IN1P[25], IN2);
  UB1BPPG_26_10 U27 (O[36], IN1P[26], IN2);
  UB1BPPG_27_10 U28 (O[37], IN1P[27], IN2);
  UB1BPPG_28_10 U29 (O[38], IN1P[28], IN2);
  UB1BPPG_29_10 U30 (O[39], IN1P[29], IN2);
  UB1BPPG_30_10 U31 (O[40], IN1P[30], IN2);
  NU1BPPG_31_10 U32 (NEG, IN1N, IN2);
  NUBUB1CON_41 U33 (O[41], NEG);
endmodule

module TCUVPPG_31_0_11 (O, IN1, IN2);
  output [42:11] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_11 U1 (O[11], IN1P[0], IN2);
  UB1BPPG_1_11 U2 (O[12], IN1P[1], IN2);
  UB1BPPG_2_11 U3 (O[13], IN1P[2], IN2);
  UB1BPPG_3_11 U4 (O[14], IN1P[3], IN2);
  UB1BPPG_4_11 U5 (O[15], IN1P[4], IN2);
  UB1BPPG_5_11 U6 (O[16], IN1P[5], IN2);
  UB1BPPG_6_11 U7 (O[17], IN1P[6], IN2);
  UB1BPPG_7_11 U8 (O[18], IN1P[7], IN2);
  UB1BPPG_8_11 U9 (O[19], IN1P[8], IN2);
  UB1BPPG_9_11 U10 (O[20], IN1P[9], IN2);
  UB1BPPG_10_11 U11 (O[21], IN1P[10], IN2);
  UB1BPPG_11_11 U12 (O[22], IN1P[11], IN2);
  UB1BPPG_12_11 U13 (O[23], IN1P[12], IN2);
  UB1BPPG_13_11 U14 (O[24], IN1P[13], IN2);
  UB1BPPG_14_11 U15 (O[25], IN1P[14], IN2);
  UB1BPPG_15_11 U16 (O[26], IN1P[15], IN2);
  UB1BPPG_16_11 U17 (O[27], IN1P[16], IN2);
  UB1BPPG_17_11 U18 (O[28], IN1P[17], IN2);
  UB1BPPG_18_11 U19 (O[29], IN1P[18], IN2);
  UB1BPPG_19_11 U20 (O[30], IN1P[19], IN2);
  UB1BPPG_20_11 U21 (O[31], IN1P[20], IN2);
  UB1BPPG_21_11 U22 (O[32], IN1P[21], IN2);
  UB1BPPG_22_11 U23 (O[33], IN1P[22], IN2);
  UB1BPPG_23_11 U24 (O[34], IN1P[23], IN2);
  UB1BPPG_24_11 U25 (O[35], IN1P[24], IN2);
  UB1BPPG_25_11 U26 (O[36], IN1P[25], IN2);
  UB1BPPG_26_11 U27 (O[37], IN1P[26], IN2);
  UB1BPPG_27_11 U28 (O[38], IN1P[27], IN2);
  UB1BPPG_28_11 U29 (O[39], IN1P[28], IN2);
  UB1BPPG_29_11 U30 (O[40], IN1P[29], IN2);
  UB1BPPG_30_11 U31 (O[41], IN1P[30], IN2);
  NU1BPPG_31_11 U32 (NEG, IN1N, IN2);
  NUBUB1CON_42 U33 (O[42], NEG);
endmodule

module TCUVPPG_31_0_12 (O, IN1, IN2);
  output [43:12] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_12 U1 (O[12], IN1P[0], IN2);
  UB1BPPG_1_12 U2 (O[13], IN1P[1], IN2);
  UB1BPPG_2_12 U3 (O[14], IN1P[2], IN2);
  UB1BPPG_3_12 U4 (O[15], IN1P[3], IN2);
  UB1BPPG_4_12 U5 (O[16], IN1P[4], IN2);
  UB1BPPG_5_12 U6 (O[17], IN1P[5], IN2);
  UB1BPPG_6_12 U7 (O[18], IN1P[6], IN2);
  UB1BPPG_7_12 U8 (O[19], IN1P[7], IN2);
  UB1BPPG_8_12 U9 (O[20], IN1P[8], IN2);
  UB1BPPG_9_12 U10 (O[21], IN1P[9], IN2);
  UB1BPPG_10_12 U11 (O[22], IN1P[10], IN2);
  UB1BPPG_11_12 U12 (O[23], IN1P[11], IN2);
  UB1BPPG_12_12 U13 (O[24], IN1P[12], IN2);
  UB1BPPG_13_12 U14 (O[25], IN1P[13], IN2);
  UB1BPPG_14_12 U15 (O[26], IN1P[14], IN2);
  UB1BPPG_15_12 U16 (O[27], IN1P[15], IN2);
  UB1BPPG_16_12 U17 (O[28], IN1P[16], IN2);
  UB1BPPG_17_12 U18 (O[29], IN1P[17], IN2);
  UB1BPPG_18_12 U19 (O[30], IN1P[18], IN2);
  UB1BPPG_19_12 U20 (O[31], IN1P[19], IN2);
  UB1BPPG_20_12 U21 (O[32], IN1P[20], IN2);
  UB1BPPG_21_12 U22 (O[33], IN1P[21], IN2);
  UB1BPPG_22_12 U23 (O[34], IN1P[22], IN2);
  UB1BPPG_23_12 U24 (O[35], IN1P[23], IN2);
  UB1BPPG_24_12 U25 (O[36], IN1P[24], IN2);
  UB1BPPG_25_12 U26 (O[37], IN1P[25], IN2);
  UB1BPPG_26_12 U27 (O[38], IN1P[26], IN2);
  UB1BPPG_27_12 U28 (O[39], IN1P[27], IN2);
  UB1BPPG_28_12 U29 (O[40], IN1P[28], IN2);
  UB1BPPG_29_12 U30 (O[41], IN1P[29], IN2);
  UB1BPPG_30_12 U31 (O[42], IN1P[30], IN2);
  NU1BPPG_31_12 U32 (NEG, IN1N, IN2);
  NUBUB1CON_43 U33 (O[43], NEG);
endmodule

module TCUVPPG_31_0_13 (O, IN1, IN2);
  output [44:13] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_13 U1 (O[13], IN1P[0], IN2);
  UB1BPPG_1_13 U2 (O[14], IN1P[1], IN2);
  UB1BPPG_2_13 U3 (O[15], IN1P[2], IN2);
  UB1BPPG_3_13 U4 (O[16], IN1P[3], IN2);
  UB1BPPG_4_13 U5 (O[17], IN1P[4], IN2);
  UB1BPPG_5_13 U6 (O[18], IN1P[5], IN2);
  UB1BPPG_6_13 U7 (O[19], IN1P[6], IN2);
  UB1BPPG_7_13 U8 (O[20], IN1P[7], IN2);
  UB1BPPG_8_13 U9 (O[21], IN1P[8], IN2);
  UB1BPPG_9_13 U10 (O[22], IN1P[9], IN2);
  UB1BPPG_10_13 U11 (O[23], IN1P[10], IN2);
  UB1BPPG_11_13 U12 (O[24], IN1P[11], IN2);
  UB1BPPG_12_13 U13 (O[25], IN1P[12], IN2);
  UB1BPPG_13_13 U14 (O[26], IN1P[13], IN2);
  UB1BPPG_14_13 U15 (O[27], IN1P[14], IN2);
  UB1BPPG_15_13 U16 (O[28], IN1P[15], IN2);
  UB1BPPG_16_13 U17 (O[29], IN1P[16], IN2);
  UB1BPPG_17_13 U18 (O[30], IN1P[17], IN2);
  UB1BPPG_18_13 U19 (O[31], IN1P[18], IN2);
  UB1BPPG_19_13 U20 (O[32], IN1P[19], IN2);
  UB1BPPG_20_13 U21 (O[33], IN1P[20], IN2);
  UB1BPPG_21_13 U22 (O[34], IN1P[21], IN2);
  UB1BPPG_22_13 U23 (O[35], IN1P[22], IN2);
  UB1BPPG_23_13 U24 (O[36], IN1P[23], IN2);
  UB1BPPG_24_13 U25 (O[37], IN1P[24], IN2);
  UB1BPPG_25_13 U26 (O[38], IN1P[25], IN2);
  UB1BPPG_26_13 U27 (O[39], IN1P[26], IN2);
  UB1BPPG_27_13 U28 (O[40], IN1P[27], IN2);
  UB1BPPG_28_13 U29 (O[41], IN1P[28], IN2);
  UB1BPPG_29_13 U30 (O[42], IN1P[29], IN2);
  UB1BPPG_30_13 U31 (O[43], IN1P[30], IN2);
  NU1BPPG_31_13 U32 (NEG, IN1N, IN2);
  NUBUB1CON_44 U33 (O[44], NEG);
endmodule

module TCUVPPG_31_0_14 (O, IN1, IN2);
  output [45:14] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_14 U1 (O[14], IN1P[0], IN2);
  UB1BPPG_1_14 U2 (O[15], IN1P[1], IN2);
  UB1BPPG_2_14 U3 (O[16], IN1P[2], IN2);
  UB1BPPG_3_14 U4 (O[17], IN1P[3], IN2);
  UB1BPPG_4_14 U5 (O[18], IN1P[4], IN2);
  UB1BPPG_5_14 U6 (O[19], IN1P[5], IN2);
  UB1BPPG_6_14 U7 (O[20], IN1P[6], IN2);
  UB1BPPG_7_14 U8 (O[21], IN1P[7], IN2);
  UB1BPPG_8_14 U9 (O[22], IN1P[8], IN2);
  UB1BPPG_9_14 U10 (O[23], IN1P[9], IN2);
  UB1BPPG_10_14 U11 (O[24], IN1P[10], IN2);
  UB1BPPG_11_14 U12 (O[25], IN1P[11], IN2);
  UB1BPPG_12_14 U13 (O[26], IN1P[12], IN2);
  UB1BPPG_13_14 U14 (O[27], IN1P[13], IN2);
  UB1BPPG_14_14 U15 (O[28], IN1P[14], IN2);
  UB1BPPG_15_14 U16 (O[29], IN1P[15], IN2);
  UB1BPPG_16_14 U17 (O[30], IN1P[16], IN2);
  UB1BPPG_17_14 U18 (O[31], IN1P[17], IN2);
  UB1BPPG_18_14 U19 (O[32], IN1P[18], IN2);
  UB1BPPG_19_14 U20 (O[33], IN1P[19], IN2);
  UB1BPPG_20_14 U21 (O[34], IN1P[20], IN2);
  UB1BPPG_21_14 U22 (O[35], IN1P[21], IN2);
  UB1BPPG_22_14 U23 (O[36], IN1P[22], IN2);
  UB1BPPG_23_14 U24 (O[37], IN1P[23], IN2);
  UB1BPPG_24_14 U25 (O[38], IN1P[24], IN2);
  UB1BPPG_25_14 U26 (O[39], IN1P[25], IN2);
  UB1BPPG_26_14 U27 (O[40], IN1P[26], IN2);
  UB1BPPG_27_14 U28 (O[41], IN1P[27], IN2);
  UB1BPPG_28_14 U29 (O[42], IN1P[28], IN2);
  UB1BPPG_29_14 U30 (O[43], IN1P[29], IN2);
  UB1BPPG_30_14 U31 (O[44], IN1P[30], IN2);
  NU1BPPG_31_14 U32 (NEG, IN1N, IN2);
  NUBUB1CON_45 U33 (O[45], NEG);
endmodule

module TCUVPPG_31_0_15 (O, IN1, IN2);
  output [46:15] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_15 U1 (O[15], IN1P[0], IN2);
  UB1BPPG_1_15 U2 (O[16], IN1P[1], IN2);
  UB1BPPG_2_15 U3 (O[17], IN1P[2], IN2);
  UB1BPPG_3_15 U4 (O[18], IN1P[3], IN2);
  UB1BPPG_4_15 U5 (O[19], IN1P[4], IN2);
  UB1BPPG_5_15 U6 (O[20], IN1P[5], IN2);
  UB1BPPG_6_15 U7 (O[21], IN1P[6], IN2);
  UB1BPPG_7_15 U8 (O[22], IN1P[7], IN2);
  UB1BPPG_8_15 U9 (O[23], IN1P[8], IN2);
  UB1BPPG_9_15 U10 (O[24], IN1P[9], IN2);
  UB1BPPG_10_15 U11 (O[25], IN1P[10], IN2);
  UB1BPPG_11_15 U12 (O[26], IN1P[11], IN2);
  UB1BPPG_12_15 U13 (O[27], IN1P[12], IN2);
  UB1BPPG_13_15 U14 (O[28], IN1P[13], IN2);
  UB1BPPG_14_15 U15 (O[29], IN1P[14], IN2);
  UB1BPPG_15_15 U16 (O[30], IN1P[15], IN2);
  UB1BPPG_16_15 U17 (O[31], IN1P[16], IN2);
  UB1BPPG_17_15 U18 (O[32], IN1P[17], IN2);
  UB1BPPG_18_15 U19 (O[33], IN1P[18], IN2);
  UB1BPPG_19_15 U20 (O[34], IN1P[19], IN2);
  UB1BPPG_20_15 U21 (O[35], IN1P[20], IN2);
  UB1BPPG_21_15 U22 (O[36], IN1P[21], IN2);
  UB1BPPG_22_15 U23 (O[37], IN1P[22], IN2);
  UB1BPPG_23_15 U24 (O[38], IN1P[23], IN2);
  UB1BPPG_24_15 U25 (O[39], IN1P[24], IN2);
  UB1BPPG_25_15 U26 (O[40], IN1P[25], IN2);
  UB1BPPG_26_15 U27 (O[41], IN1P[26], IN2);
  UB1BPPG_27_15 U28 (O[42], IN1P[27], IN2);
  UB1BPPG_28_15 U29 (O[43], IN1P[28], IN2);
  UB1BPPG_29_15 U30 (O[44], IN1P[29], IN2);
  UB1BPPG_30_15 U31 (O[45], IN1P[30], IN2);
  NU1BPPG_31_15 U32 (NEG, IN1N, IN2);
  NUBUB1CON_46 U33 (O[46], NEG);
endmodule

module TCUVPPG_31_0_16 (O, IN1, IN2);
  output [47:16] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_16 U1 (O[16], IN1P[0], IN2);
  UB1BPPG_1_16 U2 (O[17], IN1P[1], IN2);
  UB1BPPG_2_16 U3 (O[18], IN1P[2], IN2);
  UB1BPPG_3_16 U4 (O[19], IN1P[3], IN2);
  UB1BPPG_4_16 U5 (O[20], IN1P[4], IN2);
  UB1BPPG_5_16 U6 (O[21], IN1P[5], IN2);
  UB1BPPG_6_16 U7 (O[22], IN1P[6], IN2);
  UB1BPPG_7_16 U8 (O[23], IN1P[7], IN2);
  UB1BPPG_8_16 U9 (O[24], IN1P[8], IN2);
  UB1BPPG_9_16 U10 (O[25], IN1P[9], IN2);
  UB1BPPG_10_16 U11 (O[26], IN1P[10], IN2);
  UB1BPPG_11_16 U12 (O[27], IN1P[11], IN2);
  UB1BPPG_12_16 U13 (O[28], IN1P[12], IN2);
  UB1BPPG_13_16 U14 (O[29], IN1P[13], IN2);
  UB1BPPG_14_16 U15 (O[30], IN1P[14], IN2);
  UB1BPPG_15_16 U16 (O[31], IN1P[15], IN2);
  UB1BPPG_16_16 U17 (O[32], IN1P[16], IN2);
  UB1BPPG_17_16 U18 (O[33], IN1P[17], IN2);
  UB1BPPG_18_16 U19 (O[34], IN1P[18], IN2);
  UB1BPPG_19_16 U20 (O[35], IN1P[19], IN2);
  UB1BPPG_20_16 U21 (O[36], IN1P[20], IN2);
  UB1BPPG_21_16 U22 (O[37], IN1P[21], IN2);
  UB1BPPG_22_16 U23 (O[38], IN1P[22], IN2);
  UB1BPPG_23_16 U24 (O[39], IN1P[23], IN2);
  UB1BPPG_24_16 U25 (O[40], IN1P[24], IN2);
  UB1BPPG_25_16 U26 (O[41], IN1P[25], IN2);
  UB1BPPG_26_16 U27 (O[42], IN1P[26], IN2);
  UB1BPPG_27_16 U28 (O[43], IN1P[27], IN2);
  UB1BPPG_28_16 U29 (O[44], IN1P[28], IN2);
  UB1BPPG_29_16 U30 (O[45], IN1P[29], IN2);
  UB1BPPG_30_16 U31 (O[46], IN1P[30], IN2);
  NU1BPPG_31_16 U32 (NEG, IN1N, IN2);
  NUBUB1CON_47 U33 (O[47], NEG);
endmodule

module TCUVPPG_31_0_17 (O, IN1, IN2);
  output [48:17] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_17 U1 (O[17], IN1P[0], IN2);
  UB1BPPG_1_17 U2 (O[18], IN1P[1], IN2);
  UB1BPPG_2_17 U3 (O[19], IN1P[2], IN2);
  UB1BPPG_3_17 U4 (O[20], IN1P[3], IN2);
  UB1BPPG_4_17 U5 (O[21], IN1P[4], IN2);
  UB1BPPG_5_17 U6 (O[22], IN1P[5], IN2);
  UB1BPPG_6_17 U7 (O[23], IN1P[6], IN2);
  UB1BPPG_7_17 U8 (O[24], IN1P[7], IN2);
  UB1BPPG_8_17 U9 (O[25], IN1P[8], IN2);
  UB1BPPG_9_17 U10 (O[26], IN1P[9], IN2);
  UB1BPPG_10_17 U11 (O[27], IN1P[10], IN2);
  UB1BPPG_11_17 U12 (O[28], IN1P[11], IN2);
  UB1BPPG_12_17 U13 (O[29], IN1P[12], IN2);
  UB1BPPG_13_17 U14 (O[30], IN1P[13], IN2);
  UB1BPPG_14_17 U15 (O[31], IN1P[14], IN2);
  UB1BPPG_15_17 U16 (O[32], IN1P[15], IN2);
  UB1BPPG_16_17 U17 (O[33], IN1P[16], IN2);
  UB1BPPG_17_17 U18 (O[34], IN1P[17], IN2);
  UB1BPPG_18_17 U19 (O[35], IN1P[18], IN2);
  UB1BPPG_19_17 U20 (O[36], IN1P[19], IN2);
  UB1BPPG_20_17 U21 (O[37], IN1P[20], IN2);
  UB1BPPG_21_17 U22 (O[38], IN1P[21], IN2);
  UB1BPPG_22_17 U23 (O[39], IN1P[22], IN2);
  UB1BPPG_23_17 U24 (O[40], IN1P[23], IN2);
  UB1BPPG_24_17 U25 (O[41], IN1P[24], IN2);
  UB1BPPG_25_17 U26 (O[42], IN1P[25], IN2);
  UB1BPPG_26_17 U27 (O[43], IN1P[26], IN2);
  UB1BPPG_27_17 U28 (O[44], IN1P[27], IN2);
  UB1BPPG_28_17 U29 (O[45], IN1P[28], IN2);
  UB1BPPG_29_17 U30 (O[46], IN1P[29], IN2);
  UB1BPPG_30_17 U31 (O[47], IN1P[30], IN2);
  NU1BPPG_31_17 U32 (NEG, IN1N, IN2);
  NUBUB1CON_48 U33 (O[48], NEG);
endmodule

module TCUVPPG_31_0_18 (O, IN1, IN2);
  output [49:18] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_18 U1 (O[18], IN1P[0], IN2);
  UB1BPPG_1_18 U2 (O[19], IN1P[1], IN2);
  UB1BPPG_2_18 U3 (O[20], IN1P[2], IN2);
  UB1BPPG_3_18 U4 (O[21], IN1P[3], IN2);
  UB1BPPG_4_18 U5 (O[22], IN1P[4], IN2);
  UB1BPPG_5_18 U6 (O[23], IN1P[5], IN2);
  UB1BPPG_6_18 U7 (O[24], IN1P[6], IN2);
  UB1BPPG_7_18 U8 (O[25], IN1P[7], IN2);
  UB1BPPG_8_18 U9 (O[26], IN1P[8], IN2);
  UB1BPPG_9_18 U10 (O[27], IN1P[9], IN2);
  UB1BPPG_10_18 U11 (O[28], IN1P[10], IN2);
  UB1BPPG_11_18 U12 (O[29], IN1P[11], IN2);
  UB1BPPG_12_18 U13 (O[30], IN1P[12], IN2);
  UB1BPPG_13_18 U14 (O[31], IN1P[13], IN2);
  UB1BPPG_14_18 U15 (O[32], IN1P[14], IN2);
  UB1BPPG_15_18 U16 (O[33], IN1P[15], IN2);
  UB1BPPG_16_18 U17 (O[34], IN1P[16], IN2);
  UB1BPPG_17_18 U18 (O[35], IN1P[17], IN2);
  UB1BPPG_18_18 U19 (O[36], IN1P[18], IN2);
  UB1BPPG_19_18 U20 (O[37], IN1P[19], IN2);
  UB1BPPG_20_18 U21 (O[38], IN1P[20], IN2);
  UB1BPPG_21_18 U22 (O[39], IN1P[21], IN2);
  UB1BPPG_22_18 U23 (O[40], IN1P[22], IN2);
  UB1BPPG_23_18 U24 (O[41], IN1P[23], IN2);
  UB1BPPG_24_18 U25 (O[42], IN1P[24], IN2);
  UB1BPPG_25_18 U26 (O[43], IN1P[25], IN2);
  UB1BPPG_26_18 U27 (O[44], IN1P[26], IN2);
  UB1BPPG_27_18 U28 (O[45], IN1P[27], IN2);
  UB1BPPG_28_18 U29 (O[46], IN1P[28], IN2);
  UB1BPPG_29_18 U30 (O[47], IN1P[29], IN2);
  UB1BPPG_30_18 U31 (O[48], IN1P[30], IN2);
  NU1BPPG_31_18 U32 (NEG, IN1N, IN2);
  NUBUB1CON_49 U33 (O[49], NEG);
endmodule

module TCUVPPG_31_0_19 (O, IN1, IN2);
  output [50:19] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_19 U1 (O[19], IN1P[0], IN2);
  UB1BPPG_1_19 U2 (O[20], IN1P[1], IN2);
  UB1BPPG_2_19 U3 (O[21], IN1P[2], IN2);
  UB1BPPG_3_19 U4 (O[22], IN1P[3], IN2);
  UB1BPPG_4_19 U5 (O[23], IN1P[4], IN2);
  UB1BPPG_5_19 U6 (O[24], IN1P[5], IN2);
  UB1BPPG_6_19 U7 (O[25], IN1P[6], IN2);
  UB1BPPG_7_19 U8 (O[26], IN1P[7], IN2);
  UB1BPPG_8_19 U9 (O[27], IN1P[8], IN2);
  UB1BPPG_9_19 U10 (O[28], IN1P[9], IN2);
  UB1BPPG_10_19 U11 (O[29], IN1P[10], IN2);
  UB1BPPG_11_19 U12 (O[30], IN1P[11], IN2);
  UB1BPPG_12_19 U13 (O[31], IN1P[12], IN2);
  UB1BPPG_13_19 U14 (O[32], IN1P[13], IN2);
  UB1BPPG_14_19 U15 (O[33], IN1P[14], IN2);
  UB1BPPG_15_19 U16 (O[34], IN1P[15], IN2);
  UB1BPPG_16_19 U17 (O[35], IN1P[16], IN2);
  UB1BPPG_17_19 U18 (O[36], IN1P[17], IN2);
  UB1BPPG_18_19 U19 (O[37], IN1P[18], IN2);
  UB1BPPG_19_19 U20 (O[38], IN1P[19], IN2);
  UB1BPPG_20_19 U21 (O[39], IN1P[20], IN2);
  UB1BPPG_21_19 U22 (O[40], IN1P[21], IN2);
  UB1BPPG_22_19 U23 (O[41], IN1P[22], IN2);
  UB1BPPG_23_19 U24 (O[42], IN1P[23], IN2);
  UB1BPPG_24_19 U25 (O[43], IN1P[24], IN2);
  UB1BPPG_25_19 U26 (O[44], IN1P[25], IN2);
  UB1BPPG_26_19 U27 (O[45], IN1P[26], IN2);
  UB1BPPG_27_19 U28 (O[46], IN1P[27], IN2);
  UB1BPPG_28_19 U29 (O[47], IN1P[28], IN2);
  UB1BPPG_29_19 U30 (O[48], IN1P[29], IN2);
  UB1BPPG_30_19 U31 (O[49], IN1P[30], IN2);
  NU1BPPG_31_19 U32 (NEG, IN1N, IN2);
  NUBUB1CON_50 U33 (O[50], NEG);
endmodule

module TCUVPPG_31_0_2 (O, IN1, IN2);
  output [33:2] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_2 U1 (O[2], IN1P[0], IN2);
  UB1BPPG_1_2 U2 (O[3], IN1P[1], IN2);
  UB1BPPG_2_2 U3 (O[4], IN1P[2], IN2);
  UB1BPPG_3_2 U4 (O[5], IN1P[3], IN2);
  UB1BPPG_4_2 U5 (O[6], IN1P[4], IN2);
  UB1BPPG_5_2 U6 (O[7], IN1P[5], IN2);
  UB1BPPG_6_2 U7 (O[8], IN1P[6], IN2);
  UB1BPPG_7_2 U8 (O[9], IN1P[7], IN2);
  UB1BPPG_8_2 U9 (O[10], IN1P[8], IN2);
  UB1BPPG_9_2 U10 (O[11], IN1P[9], IN2);
  UB1BPPG_10_2 U11 (O[12], IN1P[10], IN2);
  UB1BPPG_11_2 U12 (O[13], IN1P[11], IN2);
  UB1BPPG_12_2 U13 (O[14], IN1P[12], IN2);
  UB1BPPG_13_2 U14 (O[15], IN1P[13], IN2);
  UB1BPPG_14_2 U15 (O[16], IN1P[14], IN2);
  UB1BPPG_15_2 U16 (O[17], IN1P[15], IN2);
  UB1BPPG_16_2 U17 (O[18], IN1P[16], IN2);
  UB1BPPG_17_2 U18 (O[19], IN1P[17], IN2);
  UB1BPPG_18_2 U19 (O[20], IN1P[18], IN2);
  UB1BPPG_19_2 U20 (O[21], IN1P[19], IN2);
  UB1BPPG_20_2 U21 (O[22], IN1P[20], IN2);
  UB1BPPG_21_2 U22 (O[23], IN1P[21], IN2);
  UB1BPPG_22_2 U23 (O[24], IN1P[22], IN2);
  UB1BPPG_23_2 U24 (O[25], IN1P[23], IN2);
  UB1BPPG_24_2 U25 (O[26], IN1P[24], IN2);
  UB1BPPG_25_2 U26 (O[27], IN1P[25], IN2);
  UB1BPPG_26_2 U27 (O[28], IN1P[26], IN2);
  UB1BPPG_27_2 U28 (O[29], IN1P[27], IN2);
  UB1BPPG_28_2 U29 (O[30], IN1P[28], IN2);
  UB1BPPG_29_2 U30 (O[31], IN1P[29], IN2);
  UB1BPPG_30_2 U31 (O[32], IN1P[30], IN2);
  NU1BPPG_31_2 U32 (NEG, IN1N, IN2);
  NUBUB1CON_33 U33 (O[33], NEG);
endmodule

module TCUVPPG_31_0_20 (O, IN1, IN2);
  output [51:20] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_20 U1 (O[20], IN1P[0], IN2);
  UB1BPPG_1_20 U2 (O[21], IN1P[1], IN2);
  UB1BPPG_2_20 U3 (O[22], IN1P[2], IN2);
  UB1BPPG_3_20 U4 (O[23], IN1P[3], IN2);
  UB1BPPG_4_20 U5 (O[24], IN1P[4], IN2);
  UB1BPPG_5_20 U6 (O[25], IN1P[5], IN2);
  UB1BPPG_6_20 U7 (O[26], IN1P[6], IN2);
  UB1BPPG_7_20 U8 (O[27], IN1P[7], IN2);
  UB1BPPG_8_20 U9 (O[28], IN1P[8], IN2);
  UB1BPPG_9_20 U10 (O[29], IN1P[9], IN2);
  UB1BPPG_10_20 U11 (O[30], IN1P[10], IN2);
  UB1BPPG_11_20 U12 (O[31], IN1P[11], IN2);
  UB1BPPG_12_20 U13 (O[32], IN1P[12], IN2);
  UB1BPPG_13_20 U14 (O[33], IN1P[13], IN2);
  UB1BPPG_14_20 U15 (O[34], IN1P[14], IN2);
  UB1BPPG_15_20 U16 (O[35], IN1P[15], IN2);
  UB1BPPG_16_20 U17 (O[36], IN1P[16], IN2);
  UB1BPPG_17_20 U18 (O[37], IN1P[17], IN2);
  UB1BPPG_18_20 U19 (O[38], IN1P[18], IN2);
  UB1BPPG_19_20 U20 (O[39], IN1P[19], IN2);
  UB1BPPG_20_20 U21 (O[40], IN1P[20], IN2);
  UB1BPPG_21_20 U22 (O[41], IN1P[21], IN2);
  UB1BPPG_22_20 U23 (O[42], IN1P[22], IN2);
  UB1BPPG_23_20 U24 (O[43], IN1P[23], IN2);
  UB1BPPG_24_20 U25 (O[44], IN1P[24], IN2);
  UB1BPPG_25_20 U26 (O[45], IN1P[25], IN2);
  UB1BPPG_26_20 U27 (O[46], IN1P[26], IN2);
  UB1BPPG_27_20 U28 (O[47], IN1P[27], IN2);
  UB1BPPG_28_20 U29 (O[48], IN1P[28], IN2);
  UB1BPPG_29_20 U30 (O[49], IN1P[29], IN2);
  UB1BPPG_30_20 U31 (O[50], IN1P[30], IN2);
  NU1BPPG_31_20 U32 (NEG, IN1N, IN2);
  NUBUB1CON_51 U33 (O[51], NEG);
endmodule

module TCUVPPG_31_0_21 (O, IN1, IN2);
  output [52:21] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_21 U1 (O[21], IN1P[0], IN2);
  UB1BPPG_1_21 U2 (O[22], IN1P[1], IN2);
  UB1BPPG_2_21 U3 (O[23], IN1P[2], IN2);
  UB1BPPG_3_21 U4 (O[24], IN1P[3], IN2);
  UB1BPPG_4_21 U5 (O[25], IN1P[4], IN2);
  UB1BPPG_5_21 U6 (O[26], IN1P[5], IN2);
  UB1BPPG_6_21 U7 (O[27], IN1P[6], IN2);
  UB1BPPG_7_21 U8 (O[28], IN1P[7], IN2);
  UB1BPPG_8_21 U9 (O[29], IN1P[8], IN2);
  UB1BPPG_9_21 U10 (O[30], IN1P[9], IN2);
  UB1BPPG_10_21 U11 (O[31], IN1P[10], IN2);
  UB1BPPG_11_21 U12 (O[32], IN1P[11], IN2);
  UB1BPPG_12_21 U13 (O[33], IN1P[12], IN2);
  UB1BPPG_13_21 U14 (O[34], IN1P[13], IN2);
  UB1BPPG_14_21 U15 (O[35], IN1P[14], IN2);
  UB1BPPG_15_21 U16 (O[36], IN1P[15], IN2);
  UB1BPPG_16_21 U17 (O[37], IN1P[16], IN2);
  UB1BPPG_17_21 U18 (O[38], IN1P[17], IN2);
  UB1BPPG_18_21 U19 (O[39], IN1P[18], IN2);
  UB1BPPG_19_21 U20 (O[40], IN1P[19], IN2);
  UB1BPPG_20_21 U21 (O[41], IN1P[20], IN2);
  UB1BPPG_21_21 U22 (O[42], IN1P[21], IN2);
  UB1BPPG_22_21 U23 (O[43], IN1P[22], IN2);
  UB1BPPG_23_21 U24 (O[44], IN1P[23], IN2);
  UB1BPPG_24_21 U25 (O[45], IN1P[24], IN2);
  UB1BPPG_25_21 U26 (O[46], IN1P[25], IN2);
  UB1BPPG_26_21 U27 (O[47], IN1P[26], IN2);
  UB1BPPG_27_21 U28 (O[48], IN1P[27], IN2);
  UB1BPPG_28_21 U29 (O[49], IN1P[28], IN2);
  UB1BPPG_29_21 U30 (O[50], IN1P[29], IN2);
  UB1BPPG_30_21 U31 (O[51], IN1P[30], IN2);
  NU1BPPG_31_21 U32 (NEG, IN1N, IN2);
  NUBUB1CON_52 U33 (O[52], NEG);
endmodule

module TCUVPPG_31_0_22 (O, IN1, IN2);
  output [53:22] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_22 U1 (O[22], IN1P[0], IN2);
  UB1BPPG_1_22 U2 (O[23], IN1P[1], IN2);
  UB1BPPG_2_22 U3 (O[24], IN1P[2], IN2);
  UB1BPPG_3_22 U4 (O[25], IN1P[3], IN2);
  UB1BPPG_4_22 U5 (O[26], IN1P[4], IN2);
  UB1BPPG_5_22 U6 (O[27], IN1P[5], IN2);
  UB1BPPG_6_22 U7 (O[28], IN1P[6], IN2);
  UB1BPPG_7_22 U8 (O[29], IN1P[7], IN2);
  UB1BPPG_8_22 U9 (O[30], IN1P[8], IN2);
  UB1BPPG_9_22 U10 (O[31], IN1P[9], IN2);
  UB1BPPG_10_22 U11 (O[32], IN1P[10], IN2);
  UB1BPPG_11_22 U12 (O[33], IN1P[11], IN2);
  UB1BPPG_12_22 U13 (O[34], IN1P[12], IN2);
  UB1BPPG_13_22 U14 (O[35], IN1P[13], IN2);
  UB1BPPG_14_22 U15 (O[36], IN1P[14], IN2);
  UB1BPPG_15_22 U16 (O[37], IN1P[15], IN2);
  UB1BPPG_16_22 U17 (O[38], IN1P[16], IN2);
  UB1BPPG_17_22 U18 (O[39], IN1P[17], IN2);
  UB1BPPG_18_22 U19 (O[40], IN1P[18], IN2);
  UB1BPPG_19_22 U20 (O[41], IN1P[19], IN2);
  UB1BPPG_20_22 U21 (O[42], IN1P[20], IN2);
  UB1BPPG_21_22 U22 (O[43], IN1P[21], IN2);
  UB1BPPG_22_22 U23 (O[44], IN1P[22], IN2);
  UB1BPPG_23_22 U24 (O[45], IN1P[23], IN2);
  UB1BPPG_24_22 U25 (O[46], IN1P[24], IN2);
  UB1BPPG_25_22 U26 (O[47], IN1P[25], IN2);
  UB1BPPG_26_22 U27 (O[48], IN1P[26], IN2);
  UB1BPPG_27_22 U28 (O[49], IN1P[27], IN2);
  UB1BPPG_28_22 U29 (O[50], IN1P[28], IN2);
  UB1BPPG_29_22 U30 (O[51], IN1P[29], IN2);
  UB1BPPG_30_22 U31 (O[52], IN1P[30], IN2);
  NU1BPPG_31_22 U32 (NEG, IN1N, IN2);
  NUBUB1CON_53 U33 (O[53], NEG);
endmodule

module TCUVPPG_31_0_23 (O, IN1, IN2);
  output [54:23] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_23 U1 (O[23], IN1P[0], IN2);
  UB1BPPG_1_23 U2 (O[24], IN1P[1], IN2);
  UB1BPPG_2_23 U3 (O[25], IN1P[2], IN2);
  UB1BPPG_3_23 U4 (O[26], IN1P[3], IN2);
  UB1BPPG_4_23 U5 (O[27], IN1P[4], IN2);
  UB1BPPG_5_23 U6 (O[28], IN1P[5], IN2);
  UB1BPPG_6_23 U7 (O[29], IN1P[6], IN2);
  UB1BPPG_7_23 U8 (O[30], IN1P[7], IN2);
  UB1BPPG_8_23 U9 (O[31], IN1P[8], IN2);
  UB1BPPG_9_23 U10 (O[32], IN1P[9], IN2);
  UB1BPPG_10_23 U11 (O[33], IN1P[10], IN2);
  UB1BPPG_11_23 U12 (O[34], IN1P[11], IN2);
  UB1BPPG_12_23 U13 (O[35], IN1P[12], IN2);
  UB1BPPG_13_23 U14 (O[36], IN1P[13], IN2);
  UB1BPPG_14_23 U15 (O[37], IN1P[14], IN2);
  UB1BPPG_15_23 U16 (O[38], IN1P[15], IN2);
  UB1BPPG_16_23 U17 (O[39], IN1P[16], IN2);
  UB1BPPG_17_23 U18 (O[40], IN1P[17], IN2);
  UB1BPPG_18_23 U19 (O[41], IN1P[18], IN2);
  UB1BPPG_19_23 U20 (O[42], IN1P[19], IN2);
  UB1BPPG_20_23 U21 (O[43], IN1P[20], IN2);
  UB1BPPG_21_23 U22 (O[44], IN1P[21], IN2);
  UB1BPPG_22_23 U23 (O[45], IN1P[22], IN2);
  UB1BPPG_23_23 U24 (O[46], IN1P[23], IN2);
  UB1BPPG_24_23 U25 (O[47], IN1P[24], IN2);
  UB1BPPG_25_23 U26 (O[48], IN1P[25], IN2);
  UB1BPPG_26_23 U27 (O[49], IN1P[26], IN2);
  UB1BPPG_27_23 U28 (O[50], IN1P[27], IN2);
  UB1BPPG_28_23 U29 (O[51], IN1P[28], IN2);
  UB1BPPG_29_23 U30 (O[52], IN1P[29], IN2);
  UB1BPPG_30_23 U31 (O[53], IN1P[30], IN2);
  NU1BPPG_31_23 U32 (NEG, IN1N, IN2);
  NUBUB1CON_54 U33 (O[54], NEG);
endmodule

module TCUVPPG_31_0_24 (O, IN1, IN2);
  output [55:24] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_24 U1 (O[24], IN1P[0], IN2);
  UB1BPPG_1_24 U2 (O[25], IN1P[1], IN2);
  UB1BPPG_2_24 U3 (O[26], IN1P[2], IN2);
  UB1BPPG_3_24 U4 (O[27], IN1P[3], IN2);
  UB1BPPG_4_24 U5 (O[28], IN1P[4], IN2);
  UB1BPPG_5_24 U6 (O[29], IN1P[5], IN2);
  UB1BPPG_6_24 U7 (O[30], IN1P[6], IN2);
  UB1BPPG_7_24 U8 (O[31], IN1P[7], IN2);
  UB1BPPG_8_24 U9 (O[32], IN1P[8], IN2);
  UB1BPPG_9_24 U10 (O[33], IN1P[9], IN2);
  UB1BPPG_10_24 U11 (O[34], IN1P[10], IN2);
  UB1BPPG_11_24 U12 (O[35], IN1P[11], IN2);
  UB1BPPG_12_24 U13 (O[36], IN1P[12], IN2);
  UB1BPPG_13_24 U14 (O[37], IN1P[13], IN2);
  UB1BPPG_14_24 U15 (O[38], IN1P[14], IN2);
  UB1BPPG_15_24 U16 (O[39], IN1P[15], IN2);
  UB1BPPG_16_24 U17 (O[40], IN1P[16], IN2);
  UB1BPPG_17_24 U18 (O[41], IN1P[17], IN2);
  UB1BPPG_18_24 U19 (O[42], IN1P[18], IN2);
  UB1BPPG_19_24 U20 (O[43], IN1P[19], IN2);
  UB1BPPG_20_24 U21 (O[44], IN1P[20], IN2);
  UB1BPPG_21_24 U22 (O[45], IN1P[21], IN2);
  UB1BPPG_22_24 U23 (O[46], IN1P[22], IN2);
  UB1BPPG_23_24 U24 (O[47], IN1P[23], IN2);
  UB1BPPG_24_24 U25 (O[48], IN1P[24], IN2);
  UB1BPPG_25_24 U26 (O[49], IN1P[25], IN2);
  UB1BPPG_26_24 U27 (O[50], IN1P[26], IN2);
  UB1BPPG_27_24 U28 (O[51], IN1P[27], IN2);
  UB1BPPG_28_24 U29 (O[52], IN1P[28], IN2);
  UB1BPPG_29_24 U30 (O[53], IN1P[29], IN2);
  UB1BPPG_30_24 U31 (O[54], IN1P[30], IN2);
  NU1BPPG_31_24 U32 (NEG, IN1N, IN2);
  NUBUB1CON_55 U33 (O[55], NEG);
endmodule

module TCUVPPG_31_0_25 (O, IN1, IN2);
  output [56:25] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_25 U1 (O[25], IN1P[0], IN2);
  UB1BPPG_1_25 U2 (O[26], IN1P[1], IN2);
  UB1BPPG_2_25 U3 (O[27], IN1P[2], IN2);
  UB1BPPG_3_25 U4 (O[28], IN1P[3], IN2);
  UB1BPPG_4_25 U5 (O[29], IN1P[4], IN2);
  UB1BPPG_5_25 U6 (O[30], IN1P[5], IN2);
  UB1BPPG_6_25 U7 (O[31], IN1P[6], IN2);
  UB1BPPG_7_25 U8 (O[32], IN1P[7], IN2);
  UB1BPPG_8_25 U9 (O[33], IN1P[8], IN2);
  UB1BPPG_9_25 U10 (O[34], IN1P[9], IN2);
  UB1BPPG_10_25 U11 (O[35], IN1P[10], IN2);
  UB1BPPG_11_25 U12 (O[36], IN1P[11], IN2);
  UB1BPPG_12_25 U13 (O[37], IN1P[12], IN2);
  UB1BPPG_13_25 U14 (O[38], IN1P[13], IN2);
  UB1BPPG_14_25 U15 (O[39], IN1P[14], IN2);
  UB1BPPG_15_25 U16 (O[40], IN1P[15], IN2);
  UB1BPPG_16_25 U17 (O[41], IN1P[16], IN2);
  UB1BPPG_17_25 U18 (O[42], IN1P[17], IN2);
  UB1BPPG_18_25 U19 (O[43], IN1P[18], IN2);
  UB1BPPG_19_25 U20 (O[44], IN1P[19], IN2);
  UB1BPPG_20_25 U21 (O[45], IN1P[20], IN2);
  UB1BPPG_21_25 U22 (O[46], IN1P[21], IN2);
  UB1BPPG_22_25 U23 (O[47], IN1P[22], IN2);
  UB1BPPG_23_25 U24 (O[48], IN1P[23], IN2);
  UB1BPPG_24_25 U25 (O[49], IN1P[24], IN2);
  UB1BPPG_25_25 U26 (O[50], IN1P[25], IN2);
  UB1BPPG_26_25 U27 (O[51], IN1P[26], IN2);
  UB1BPPG_27_25 U28 (O[52], IN1P[27], IN2);
  UB1BPPG_28_25 U29 (O[53], IN1P[28], IN2);
  UB1BPPG_29_25 U30 (O[54], IN1P[29], IN2);
  UB1BPPG_30_25 U31 (O[55], IN1P[30], IN2);
  NU1BPPG_31_25 U32 (NEG, IN1N, IN2);
  NUBUB1CON_56 U33 (O[56], NEG);
endmodule

module TCUVPPG_31_0_26 (O, IN1, IN2);
  output [57:26] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_26 U1 (O[26], IN1P[0], IN2);
  UB1BPPG_1_26 U2 (O[27], IN1P[1], IN2);
  UB1BPPG_2_26 U3 (O[28], IN1P[2], IN2);
  UB1BPPG_3_26 U4 (O[29], IN1P[3], IN2);
  UB1BPPG_4_26 U5 (O[30], IN1P[4], IN2);
  UB1BPPG_5_26 U6 (O[31], IN1P[5], IN2);
  UB1BPPG_6_26 U7 (O[32], IN1P[6], IN2);
  UB1BPPG_7_26 U8 (O[33], IN1P[7], IN2);
  UB1BPPG_8_26 U9 (O[34], IN1P[8], IN2);
  UB1BPPG_9_26 U10 (O[35], IN1P[9], IN2);
  UB1BPPG_10_26 U11 (O[36], IN1P[10], IN2);
  UB1BPPG_11_26 U12 (O[37], IN1P[11], IN2);
  UB1BPPG_12_26 U13 (O[38], IN1P[12], IN2);
  UB1BPPG_13_26 U14 (O[39], IN1P[13], IN2);
  UB1BPPG_14_26 U15 (O[40], IN1P[14], IN2);
  UB1BPPG_15_26 U16 (O[41], IN1P[15], IN2);
  UB1BPPG_16_26 U17 (O[42], IN1P[16], IN2);
  UB1BPPG_17_26 U18 (O[43], IN1P[17], IN2);
  UB1BPPG_18_26 U19 (O[44], IN1P[18], IN2);
  UB1BPPG_19_26 U20 (O[45], IN1P[19], IN2);
  UB1BPPG_20_26 U21 (O[46], IN1P[20], IN2);
  UB1BPPG_21_26 U22 (O[47], IN1P[21], IN2);
  UB1BPPG_22_26 U23 (O[48], IN1P[22], IN2);
  UB1BPPG_23_26 U24 (O[49], IN1P[23], IN2);
  UB1BPPG_24_26 U25 (O[50], IN1P[24], IN2);
  UB1BPPG_25_26 U26 (O[51], IN1P[25], IN2);
  UB1BPPG_26_26 U27 (O[52], IN1P[26], IN2);
  UB1BPPG_27_26 U28 (O[53], IN1P[27], IN2);
  UB1BPPG_28_26 U29 (O[54], IN1P[28], IN2);
  UB1BPPG_29_26 U30 (O[55], IN1P[29], IN2);
  UB1BPPG_30_26 U31 (O[56], IN1P[30], IN2);
  NU1BPPG_31_26 U32 (NEG, IN1N, IN2);
  NUBUB1CON_57 U33 (O[57], NEG);
endmodule

module TCUVPPG_31_0_27 (O, IN1, IN2);
  output [58:27] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_27 U1 (O[27], IN1P[0], IN2);
  UB1BPPG_1_27 U2 (O[28], IN1P[1], IN2);
  UB1BPPG_2_27 U3 (O[29], IN1P[2], IN2);
  UB1BPPG_3_27 U4 (O[30], IN1P[3], IN2);
  UB1BPPG_4_27 U5 (O[31], IN1P[4], IN2);
  UB1BPPG_5_27 U6 (O[32], IN1P[5], IN2);
  UB1BPPG_6_27 U7 (O[33], IN1P[6], IN2);
  UB1BPPG_7_27 U8 (O[34], IN1P[7], IN2);
  UB1BPPG_8_27 U9 (O[35], IN1P[8], IN2);
  UB1BPPG_9_27 U10 (O[36], IN1P[9], IN2);
  UB1BPPG_10_27 U11 (O[37], IN1P[10], IN2);
  UB1BPPG_11_27 U12 (O[38], IN1P[11], IN2);
  UB1BPPG_12_27 U13 (O[39], IN1P[12], IN2);
  UB1BPPG_13_27 U14 (O[40], IN1P[13], IN2);
  UB1BPPG_14_27 U15 (O[41], IN1P[14], IN2);
  UB1BPPG_15_27 U16 (O[42], IN1P[15], IN2);
  UB1BPPG_16_27 U17 (O[43], IN1P[16], IN2);
  UB1BPPG_17_27 U18 (O[44], IN1P[17], IN2);
  UB1BPPG_18_27 U19 (O[45], IN1P[18], IN2);
  UB1BPPG_19_27 U20 (O[46], IN1P[19], IN2);
  UB1BPPG_20_27 U21 (O[47], IN1P[20], IN2);
  UB1BPPG_21_27 U22 (O[48], IN1P[21], IN2);
  UB1BPPG_22_27 U23 (O[49], IN1P[22], IN2);
  UB1BPPG_23_27 U24 (O[50], IN1P[23], IN2);
  UB1BPPG_24_27 U25 (O[51], IN1P[24], IN2);
  UB1BPPG_25_27 U26 (O[52], IN1P[25], IN2);
  UB1BPPG_26_27 U27 (O[53], IN1P[26], IN2);
  UB1BPPG_27_27 U28 (O[54], IN1P[27], IN2);
  UB1BPPG_28_27 U29 (O[55], IN1P[28], IN2);
  UB1BPPG_29_27 U30 (O[56], IN1P[29], IN2);
  UB1BPPG_30_27 U31 (O[57], IN1P[30], IN2);
  NU1BPPG_31_27 U32 (NEG, IN1N, IN2);
  NUBUB1CON_58 U33 (O[58], NEG);
endmodule

module TCUVPPG_31_0_28 (O, IN1, IN2);
  output [59:28] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_28 U1 (O[28], IN1P[0], IN2);
  UB1BPPG_1_28 U2 (O[29], IN1P[1], IN2);
  UB1BPPG_2_28 U3 (O[30], IN1P[2], IN2);
  UB1BPPG_3_28 U4 (O[31], IN1P[3], IN2);
  UB1BPPG_4_28 U5 (O[32], IN1P[4], IN2);
  UB1BPPG_5_28 U6 (O[33], IN1P[5], IN2);
  UB1BPPG_6_28 U7 (O[34], IN1P[6], IN2);
  UB1BPPG_7_28 U8 (O[35], IN1P[7], IN2);
  UB1BPPG_8_28 U9 (O[36], IN1P[8], IN2);
  UB1BPPG_9_28 U10 (O[37], IN1P[9], IN2);
  UB1BPPG_10_28 U11 (O[38], IN1P[10], IN2);
  UB1BPPG_11_28 U12 (O[39], IN1P[11], IN2);
  UB1BPPG_12_28 U13 (O[40], IN1P[12], IN2);
  UB1BPPG_13_28 U14 (O[41], IN1P[13], IN2);
  UB1BPPG_14_28 U15 (O[42], IN1P[14], IN2);
  UB1BPPG_15_28 U16 (O[43], IN1P[15], IN2);
  UB1BPPG_16_28 U17 (O[44], IN1P[16], IN2);
  UB1BPPG_17_28 U18 (O[45], IN1P[17], IN2);
  UB1BPPG_18_28 U19 (O[46], IN1P[18], IN2);
  UB1BPPG_19_28 U20 (O[47], IN1P[19], IN2);
  UB1BPPG_20_28 U21 (O[48], IN1P[20], IN2);
  UB1BPPG_21_28 U22 (O[49], IN1P[21], IN2);
  UB1BPPG_22_28 U23 (O[50], IN1P[22], IN2);
  UB1BPPG_23_28 U24 (O[51], IN1P[23], IN2);
  UB1BPPG_24_28 U25 (O[52], IN1P[24], IN2);
  UB1BPPG_25_28 U26 (O[53], IN1P[25], IN2);
  UB1BPPG_26_28 U27 (O[54], IN1P[26], IN2);
  UB1BPPG_27_28 U28 (O[55], IN1P[27], IN2);
  UB1BPPG_28_28 U29 (O[56], IN1P[28], IN2);
  UB1BPPG_29_28 U30 (O[57], IN1P[29], IN2);
  UB1BPPG_30_28 U31 (O[58], IN1P[30], IN2);
  NU1BPPG_31_28 U32 (NEG, IN1N, IN2);
  NUBUB1CON_59 U33 (O[59], NEG);
endmodule

module TCUVPPG_31_0_29 (O, IN1, IN2);
  output [60:29] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_29 U1 (O[29], IN1P[0], IN2);
  UB1BPPG_1_29 U2 (O[30], IN1P[1], IN2);
  UB1BPPG_2_29 U3 (O[31], IN1P[2], IN2);
  UB1BPPG_3_29 U4 (O[32], IN1P[3], IN2);
  UB1BPPG_4_29 U5 (O[33], IN1P[4], IN2);
  UB1BPPG_5_29 U6 (O[34], IN1P[5], IN2);
  UB1BPPG_6_29 U7 (O[35], IN1P[6], IN2);
  UB1BPPG_7_29 U8 (O[36], IN1P[7], IN2);
  UB1BPPG_8_29 U9 (O[37], IN1P[8], IN2);
  UB1BPPG_9_29 U10 (O[38], IN1P[9], IN2);
  UB1BPPG_10_29 U11 (O[39], IN1P[10], IN2);
  UB1BPPG_11_29 U12 (O[40], IN1P[11], IN2);
  UB1BPPG_12_29 U13 (O[41], IN1P[12], IN2);
  UB1BPPG_13_29 U14 (O[42], IN1P[13], IN2);
  UB1BPPG_14_29 U15 (O[43], IN1P[14], IN2);
  UB1BPPG_15_29 U16 (O[44], IN1P[15], IN2);
  UB1BPPG_16_29 U17 (O[45], IN1P[16], IN2);
  UB1BPPG_17_29 U18 (O[46], IN1P[17], IN2);
  UB1BPPG_18_29 U19 (O[47], IN1P[18], IN2);
  UB1BPPG_19_29 U20 (O[48], IN1P[19], IN2);
  UB1BPPG_20_29 U21 (O[49], IN1P[20], IN2);
  UB1BPPG_21_29 U22 (O[50], IN1P[21], IN2);
  UB1BPPG_22_29 U23 (O[51], IN1P[22], IN2);
  UB1BPPG_23_29 U24 (O[52], IN1P[23], IN2);
  UB1BPPG_24_29 U25 (O[53], IN1P[24], IN2);
  UB1BPPG_25_29 U26 (O[54], IN1P[25], IN2);
  UB1BPPG_26_29 U27 (O[55], IN1P[26], IN2);
  UB1BPPG_27_29 U28 (O[56], IN1P[27], IN2);
  UB1BPPG_28_29 U29 (O[57], IN1P[28], IN2);
  UB1BPPG_29_29 U30 (O[58], IN1P[29], IN2);
  UB1BPPG_30_29 U31 (O[59], IN1P[30], IN2);
  NU1BPPG_31_29 U32 (NEG, IN1N, IN2);
  NUBUB1CON_60 U33 (O[60], NEG);
endmodule

module TCUVPPG_31_0_3 (O, IN1, IN2);
  output [34:3] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_3 U1 (O[3], IN1P[0], IN2);
  UB1BPPG_1_3 U2 (O[4], IN1P[1], IN2);
  UB1BPPG_2_3 U3 (O[5], IN1P[2], IN2);
  UB1BPPG_3_3 U4 (O[6], IN1P[3], IN2);
  UB1BPPG_4_3 U5 (O[7], IN1P[4], IN2);
  UB1BPPG_5_3 U6 (O[8], IN1P[5], IN2);
  UB1BPPG_6_3 U7 (O[9], IN1P[6], IN2);
  UB1BPPG_7_3 U8 (O[10], IN1P[7], IN2);
  UB1BPPG_8_3 U9 (O[11], IN1P[8], IN2);
  UB1BPPG_9_3 U10 (O[12], IN1P[9], IN2);
  UB1BPPG_10_3 U11 (O[13], IN1P[10], IN2);
  UB1BPPG_11_3 U12 (O[14], IN1P[11], IN2);
  UB1BPPG_12_3 U13 (O[15], IN1P[12], IN2);
  UB1BPPG_13_3 U14 (O[16], IN1P[13], IN2);
  UB1BPPG_14_3 U15 (O[17], IN1P[14], IN2);
  UB1BPPG_15_3 U16 (O[18], IN1P[15], IN2);
  UB1BPPG_16_3 U17 (O[19], IN1P[16], IN2);
  UB1BPPG_17_3 U18 (O[20], IN1P[17], IN2);
  UB1BPPG_18_3 U19 (O[21], IN1P[18], IN2);
  UB1BPPG_19_3 U20 (O[22], IN1P[19], IN2);
  UB1BPPG_20_3 U21 (O[23], IN1P[20], IN2);
  UB1BPPG_21_3 U22 (O[24], IN1P[21], IN2);
  UB1BPPG_22_3 U23 (O[25], IN1P[22], IN2);
  UB1BPPG_23_3 U24 (O[26], IN1P[23], IN2);
  UB1BPPG_24_3 U25 (O[27], IN1P[24], IN2);
  UB1BPPG_25_3 U26 (O[28], IN1P[25], IN2);
  UB1BPPG_26_3 U27 (O[29], IN1P[26], IN2);
  UB1BPPG_27_3 U28 (O[30], IN1P[27], IN2);
  UB1BPPG_28_3 U29 (O[31], IN1P[28], IN2);
  UB1BPPG_29_3 U30 (O[32], IN1P[29], IN2);
  UB1BPPG_30_3 U31 (O[33], IN1P[30], IN2);
  NU1BPPG_31_3 U32 (NEG, IN1N, IN2);
  NUBUB1CON_34 U33 (O[34], NEG);
endmodule

module TCUVPPG_31_0_30 (O, IN1, IN2);
  output [61:30] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_30 U1 (O[30], IN1P[0], IN2);
  UB1BPPG_1_30 U2 (O[31], IN1P[1], IN2);
  UB1BPPG_2_30 U3 (O[32], IN1P[2], IN2);
  UB1BPPG_3_30 U4 (O[33], IN1P[3], IN2);
  UB1BPPG_4_30 U5 (O[34], IN1P[4], IN2);
  UB1BPPG_5_30 U6 (O[35], IN1P[5], IN2);
  UB1BPPG_6_30 U7 (O[36], IN1P[6], IN2);
  UB1BPPG_7_30 U8 (O[37], IN1P[7], IN2);
  UB1BPPG_8_30 U9 (O[38], IN1P[8], IN2);
  UB1BPPG_9_30 U10 (O[39], IN1P[9], IN2);
  UB1BPPG_10_30 U11 (O[40], IN1P[10], IN2);
  UB1BPPG_11_30 U12 (O[41], IN1P[11], IN2);
  UB1BPPG_12_30 U13 (O[42], IN1P[12], IN2);
  UB1BPPG_13_30 U14 (O[43], IN1P[13], IN2);
  UB1BPPG_14_30 U15 (O[44], IN1P[14], IN2);
  UB1BPPG_15_30 U16 (O[45], IN1P[15], IN2);
  UB1BPPG_16_30 U17 (O[46], IN1P[16], IN2);
  UB1BPPG_17_30 U18 (O[47], IN1P[17], IN2);
  UB1BPPG_18_30 U19 (O[48], IN1P[18], IN2);
  UB1BPPG_19_30 U20 (O[49], IN1P[19], IN2);
  UB1BPPG_20_30 U21 (O[50], IN1P[20], IN2);
  UB1BPPG_21_30 U22 (O[51], IN1P[21], IN2);
  UB1BPPG_22_30 U23 (O[52], IN1P[22], IN2);
  UB1BPPG_23_30 U24 (O[53], IN1P[23], IN2);
  UB1BPPG_24_30 U25 (O[54], IN1P[24], IN2);
  UB1BPPG_25_30 U26 (O[55], IN1P[25], IN2);
  UB1BPPG_26_30 U27 (O[56], IN1P[26], IN2);
  UB1BPPG_27_30 U28 (O[57], IN1P[27], IN2);
  UB1BPPG_28_30 U29 (O[58], IN1P[28], IN2);
  UB1BPPG_29_30 U30 (O[59], IN1P[29], IN2);
  UB1BPPG_30_30 U31 (O[60], IN1P[30], IN2);
  NU1BPPG_31_30 U32 (NEG, IN1N, IN2);
  NUBUB1CON_61 U33 (O[61], NEG);
endmodule

module TCUVPPG_31_0_4 (O, IN1, IN2);
  output [35:4] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_4 U1 (O[4], IN1P[0], IN2);
  UB1BPPG_1_4 U2 (O[5], IN1P[1], IN2);
  UB1BPPG_2_4 U3 (O[6], IN1P[2], IN2);
  UB1BPPG_3_4 U4 (O[7], IN1P[3], IN2);
  UB1BPPG_4_4 U5 (O[8], IN1P[4], IN2);
  UB1BPPG_5_4 U6 (O[9], IN1P[5], IN2);
  UB1BPPG_6_4 U7 (O[10], IN1P[6], IN2);
  UB1BPPG_7_4 U8 (O[11], IN1P[7], IN2);
  UB1BPPG_8_4 U9 (O[12], IN1P[8], IN2);
  UB1BPPG_9_4 U10 (O[13], IN1P[9], IN2);
  UB1BPPG_10_4 U11 (O[14], IN1P[10], IN2);
  UB1BPPG_11_4 U12 (O[15], IN1P[11], IN2);
  UB1BPPG_12_4 U13 (O[16], IN1P[12], IN2);
  UB1BPPG_13_4 U14 (O[17], IN1P[13], IN2);
  UB1BPPG_14_4 U15 (O[18], IN1P[14], IN2);
  UB1BPPG_15_4 U16 (O[19], IN1P[15], IN2);
  UB1BPPG_16_4 U17 (O[20], IN1P[16], IN2);
  UB1BPPG_17_4 U18 (O[21], IN1P[17], IN2);
  UB1BPPG_18_4 U19 (O[22], IN1P[18], IN2);
  UB1BPPG_19_4 U20 (O[23], IN1P[19], IN2);
  UB1BPPG_20_4 U21 (O[24], IN1P[20], IN2);
  UB1BPPG_21_4 U22 (O[25], IN1P[21], IN2);
  UB1BPPG_22_4 U23 (O[26], IN1P[22], IN2);
  UB1BPPG_23_4 U24 (O[27], IN1P[23], IN2);
  UB1BPPG_24_4 U25 (O[28], IN1P[24], IN2);
  UB1BPPG_25_4 U26 (O[29], IN1P[25], IN2);
  UB1BPPG_26_4 U27 (O[30], IN1P[26], IN2);
  UB1BPPG_27_4 U28 (O[31], IN1P[27], IN2);
  UB1BPPG_28_4 U29 (O[32], IN1P[28], IN2);
  UB1BPPG_29_4 U30 (O[33], IN1P[29], IN2);
  UB1BPPG_30_4 U31 (O[34], IN1P[30], IN2);
  NU1BPPG_31_4 U32 (NEG, IN1N, IN2);
  NUBUB1CON_35 U33 (O[35], NEG);
endmodule

module TCUVPPG_31_0_5 (O, IN1, IN2);
  output [36:5] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_5 U1 (O[5], IN1P[0], IN2);
  UB1BPPG_1_5 U2 (O[6], IN1P[1], IN2);
  UB1BPPG_2_5 U3 (O[7], IN1P[2], IN2);
  UB1BPPG_3_5 U4 (O[8], IN1P[3], IN2);
  UB1BPPG_4_5 U5 (O[9], IN1P[4], IN2);
  UB1BPPG_5_5 U6 (O[10], IN1P[5], IN2);
  UB1BPPG_6_5 U7 (O[11], IN1P[6], IN2);
  UB1BPPG_7_5 U8 (O[12], IN1P[7], IN2);
  UB1BPPG_8_5 U9 (O[13], IN1P[8], IN2);
  UB1BPPG_9_5 U10 (O[14], IN1P[9], IN2);
  UB1BPPG_10_5 U11 (O[15], IN1P[10], IN2);
  UB1BPPG_11_5 U12 (O[16], IN1P[11], IN2);
  UB1BPPG_12_5 U13 (O[17], IN1P[12], IN2);
  UB1BPPG_13_5 U14 (O[18], IN1P[13], IN2);
  UB1BPPG_14_5 U15 (O[19], IN1P[14], IN2);
  UB1BPPG_15_5 U16 (O[20], IN1P[15], IN2);
  UB1BPPG_16_5 U17 (O[21], IN1P[16], IN2);
  UB1BPPG_17_5 U18 (O[22], IN1P[17], IN2);
  UB1BPPG_18_5 U19 (O[23], IN1P[18], IN2);
  UB1BPPG_19_5 U20 (O[24], IN1P[19], IN2);
  UB1BPPG_20_5 U21 (O[25], IN1P[20], IN2);
  UB1BPPG_21_5 U22 (O[26], IN1P[21], IN2);
  UB1BPPG_22_5 U23 (O[27], IN1P[22], IN2);
  UB1BPPG_23_5 U24 (O[28], IN1P[23], IN2);
  UB1BPPG_24_5 U25 (O[29], IN1P[24], IN2);
  UB1BPPG_25_5 U26 (O[30], IN1P[25], IN2);
  UB1BPPG_26_5 U27 (O[31], IN1P[26], IN2);
  UB1BPPG_27_5 U28 (O[32], IN1P[27], IN2);
  UB1BPPG_28_5 U29 (O[33], IN1P[28], IN2);
  UB1BPPG_29_5 U30 (O[34], IN1P[29], IN2);
  UB1BPPG_30_5 U31 (O[35], IN1P[30], IN2);
  NU1BPPG_31_5 U32 (NEG, IN1N, IN2);
  NUBUB1CON_36 U33 (O[36], NEG);
endmodule

module TCUVPPG_31_0_6 (O, IN1, IN2);
  output [37:6] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_6 U1 (O[6], IN1P[0], IN2);
  UB1BPPG_1_6 U2 (O[7], IN1P[1], IN2);
  UB1BPPG_2_6 U3 (O[8], IN1P[2], IN2);
  UB1BPPG_3_6 U4 (O[9], IN1P[3], IN2);
  UB1BPPG_4_6 U5 (O[10], IN1P[4], IN2);
  UB1BPPG_5_6 U6 (O[11], IN1P[5], IN2);
  UB1BPPG_6_6 U7 (O[12], IN1P[6], IN2);
  UB1BPPG_7_6 U8 (O[13], IN1P[7], IN2);
  UB1BPPG_8_6 U9 (O[14], IN1P[8], IN2);
  UB1BPPG_9_6 U10 (O[15], IN1P[9], IN2);
  UB1BPPG_10_6 U11 (O[16], IN1P[10], IN2);
  UB1BPPG_11_6 U12 (O[17], IN1P[11], IN2);
  UB1BPPG_12_6 U13 (O[18], IN1P[12], IN2);
  UB1BPPG_13_6 U14 (O[19], IN1P[13], IN2);
  UB1BPPG_14_6 U15 (O[20], IN1P[14], IN2);
  UB1BPPG_15_6 U16 (O[21], IN1P[15], IN2);
  UB1BPPG_16_6 U17 (O[22], IN1P[16], IN2);
  UB1BPPG_17_6 U18 (O[23], IN1P[17], IN2);
  UB1BPPG_18_6 U19 (O[24], IN1P[18], IN2);
  UB1BPPG_19_6 U20 (O[25], IN1P[19], IN2);
  UB1BPPG_20_6 U21 (O[26], IN1P[20], IN2);
  UB1BPPG_21_6 U22 (O[27], IN1P[21], IN2);
  UB1BPPG_22_6 U23 (O[28], IN1P[22], IN2);
  UB1BPPG_23_6 U24 (O[29], IN1P[23], IN2);
  UB1BPPG_24_6 U25 (O[30], IN1P[24], IN2);
  UB1BPPG_25_6 U26 (O[31], IN1P[25], IN2);
  UB1BPPG_26_6 U27 (O[32], IN1P[26], IN2);
  UB1BPPG_27_6 U28 (O[33], IN1P[27], IN2);
  UB1BPPG_28_6 U29 (O[34], IN1P[28], IN2);
  UB1BPPG_29_6 U30 (O[35], IN1P[29], IN2);
  UB1BPPG_30_6 U31 (O[36], IN1P[30], IN2);
  NU1BPPG_31_6 U32 (NEG, IN1N, IN2);
  NUBUB1CON_37 U33 (O[37], NEG);
endmodule

module TCUVPPG_31_0_7 (O, IN1, IN2);
  output [38:7] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_7 U1 (O[7], IN1P[0], IN2);
  UB1BPPG_1_7 U2 (O[8], IN1P[1], IN2);
  UB1BPPG_2_7 U3 (O[9], IN1P[2], IN2);
  UB1BPPG_3_7 U4 (O[10], IN1P[3], IN2);
  UB1BPPG_4_7 U5 (O[11], IN1P[4], IN2);
  UB1BPPG_5_7 U6 (O[12], IN1P[5], IN2);
  UB1BPPG_6_7 U7 (O[13], IN1P[6], IN2);
  UB1BPPG_7_7 U8 (O[14], IN1P[7], IN2);
  UB1BPPG_8_7 U9 (O[15], IN1P[8], IN2);
  UB1BPPG_9_7 U10 (O[16], IN1P[9], IN2);
  UB1BPPG_10_7 U11 (O[17], IN1P[10], IN2);
  UB1BPPG_11_7 U12 (O[18], IN1P[11], IN2);
  UB1BPPG_12_7 U13 (O[19], IN1P[12], IN2);
  UB1BPPG_13_7 U14 (O[20], IN1P[13], IN2);
  UB1BPPG_14_7 U15 (O[21], IN1P[14], IN2);
  UB1BPPG_15_7 U16 (O[22], IN1P[15], IN2);
  UB1BPPG_16_7 U17 (O[23], IN1P[16], IN2);
  UB1BPPG_17_7 U18 (O[24], IN1P[17], IN2);
  UB1BPPG_18_7 U19 (O[25], IN1P[18], IN2);
  UB1BPPG_19_7 U20 (O[26], IN1P[19], IN2);
  UB1BPPG_20_7 U21 (O[27], IN1P[20], IN2);
  UB1BPPG_21_7 U22 (O[28], IN1P[21], IN2);
  UB1BPPG_22_7 U23 (O[29], IN1P[22], IN2);
  UB1BPPG_23_7 U24 (O[30], IN1P[23], IN2);
  UB1BPPG_24_7 U25 (O[31], IN1P[24], IN2);
  UB1BPPG_25_7 U26 (O[32], IN1P[25], IN2);
  UB1BPPG_26_7 U27 (O[33], IN1P[26], IN2);
  UB1BPPG_27_7 U28 (O[34], IN1P[27], IN2);
  UB1BPPG_28_7 U29 (O[35], IN1P[28], IN2);
  UB1BPPG_29_7 U30 (O[36], IN1P[29], IN2);
  UB1BPPG_30_7 U31 (O[37], IN1P[30], IN2);
  NU1BPPG_31_7 U32 (NEG, IN1N, IN2);
  NUBUB1CON_38 U33 (O[38], NEG);
endmodule

module TCUVPPG_31_0_8 (O, IN1, IN2);
  output [39:8] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_8 U1 (O[8], IN1P[0], IN2);
  UB1BPPG_1_8 U2 (O[9], IN1P[1], IN2);
  UB1BPPG_2_8 U3 (O[10], IN1P[2], IN2);
  UB1BPPG_3_8 U4 (O[11], IN1P[3], IN2);
  UB1BPPG_4_8 U5 (O[12], IN1P[4], IN2);
  UB1BPPG_5_8 U6 (O[13], IN1P[5], IN2);
  UB1BPPG_6_8 U7 (O[14], IN1P[6], IN2);
  UB1BPPG_7_8 U8 (O[15], IN1P[7], IN2);
  UB1BPPG_8_8 U9 (O[16], IN1P[8], IN2);
  UB1BPPG_9_8 U10 (O[17], IN1P[9], IN2);
  UB1BPPG_10_8 U11 (O[18], IN1P[10], IN2);
  UB1BPPG_11_8 U12 (O[19], IN1P[11], IN2);
  UB1BPPG_12_8 U13 (O[20], IN1P[12], IN2);
  UB1BPPG_13_8 U14 (O[21], IN1P[13], IN2);
  UB1BPPG_14_8 U15 (O[22], IN1P[14], IN2);
  UB1BPPG_15_8 U16 (O[23], IN1P[15], IN2);
  UB1BPPG_16_8 U17 (O[24], IN1P[16], IN2);
  UB1BPPG_17_8 U18 (O[25], IN1P[17], IN2);
  UB1BPPG_18_8 U19 (O[26], IN1P[18], IN2);
  UB1BPPG_19_8 U20 (O[27], IN1P[19], IN2);
  UB1BPPG_20_8 U21 (O[28], IN1P[20], IN2);
  UB1BPPG_21_8 U22 (O[29], IN1P[21], IN2);
  UB1BPPG_22_8 U23 (O[30], IN1P[22], IN2);
  UB1BPPG_23_8 U24 (O[31], IN1P[23], IN2);
  UB1BPPG_24_8 U25 (O[32], IN1P[24], IN2);
  UB1BPPG_25_8 U26 (O[33], IN1P[25], IN2);
  UB1BPPG_26_8 U27 (O[34], IN1P[26], IN2);
  UB1BPPG_27_8 U28 (O[35], IN1P[27], IN2);
  UB1BPPG_28_8 U29 (O[36], IN1P[28], IN2);
  UB1BPPG_29_8 U30 (O[37], IN1P[29], IN2);
  UB1BPPG_30_8 U31 (O[38], IN1P[30], IN2);
  NU1BPPG_31_8 U32 (NEG, IN1N, IN2);
  NUBUB1CON_39 U33 (O[39], NEG);
endmodule

module TCUVPPG_31_0_9 (O, IN1, IN2);
  output [40:9] O;
  input [31:0] IN1;
  input IN2;
  wire IN1N;
  wire [30:0] IN1P;
  wire NEG;
  TCDECON_31_0 U0 (IN1N, IN1P, IN1);
  UB1BPPG_0_9 U1 (O[9], IN1P[0], IN2);
  UB1BPPG_1_9 U2 (O[10], IN1P[1], IN2);
  UB1BPPG_2_9 U3 (O[11], IN1P[2], IN2);
  UB1BPPG_3_9 U4 (O[12], IN1P[3], IN2);
  UB1BPPG_4_9 U5 (O[13], IN1P[4], IN2);
  UB1BPPG_5_9 U6 (O[14], IN1P[5], IN2);
  UB1BPPG_6_9 U7 (O[15], IN1P[6], IN2);
  UB1BPPG_7_9 U8 (O[16], IN1P[7], IN2);
  UB1BPPG_8_9 U9 (O[17], IN1P[8], IN2);
  UB1BPPG_9_9 U10 (O[18], IN1P[9], IN2);
  UB1BPPG_10_9 U11 (O[19], IN1P[10], IN2);
  UB1BPPG_11_9 U12 (O[20], IN1P[11], IN2);
  UB1BPPG_12_9 U13 (O[21], IN1P[12], IN2);
  UB1BPPG_13_9 U14 (O[22], IN1P[13], IN2);
  UB1BPPG_14_9 U15 (O[23], IN1P[14], IN2);
  UB1BPPG_15_9 U16 (O[24], IN1P[15], IN2);
  UB1BPPG_16_9 U17 (O[25], IN1P[16], IN2);
  UB1BPPG_17_9 U18 (O[26], IN1P[17], IN2);
  UB1BPPG_18_9 U19 (O[27], IN1P[18], IN2);
  UB1BPPG_19_9 U20 (O[28], IN1P[19], IN2);
  UB1BPPG_20_9 U21 (O[29], IN1P[20], IN2);
  UB1BPPG_21_9 U22 (O[30], IN1P[21], IN2);
  UB1BPPG_22_9 U23 (O[31], IN1P[22], IN2);
  UB1BPPG_23_9 U24 (O[32], IN1P[23], IN2);
  UB1BPPG_24_9 U25 (O[33], IN1P[24], IN2);
  UB1BPPG_25_9 U26 (O[34], IN1P[25], IN2);
  UB1BPPG_26_9 U27 (O[35], IN1P[26], IN2);
  UB1BPPG_27_9 U28 (O[36], IN1P[27], IN2);
  UB1BPPG_28_9 U29 (O[37], IN1P[28], IN2);
  UB1BPPG_29_9 U30 (O[38], IN1P[29], IN2);
  UB1BPPG_30_9 U31 (O[39], IN1P[30], IN2);
  NU1BPPG_31_9 U32 (NEG, IN1N, IN2);
  NUBUB1CON_40 U33 (O[40], NEG);
endmodule

module UBCMBIN_32_32_31_000 (O, IN0, IN1);
  output [32:0] O;
  input IN0;
  input [31:0] IN1;
  UB1DCON_32 U0 (O[32], IN0);
  UBCON_31_0 U1 (O[31:0], IN1);
endmodule

module UBCON_10_9 (O, I);
  output [10:9] O;
  input [10:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
endmodule

module UBCON_12_10 (O, I);
  output [12:10] O;
  input [12:10] I;
  UB1DCON_10 U0 (O[10], I[10]);
  UB1DCON_11 U1 (O[11], I[11]);
  UB1DCON_12 U2 (O[12], I[12]);
endmodule

module UBCON_14_13 (O, I);
  output [14:13] O;
  input [14:13] I;
  UB1DCON_13 U0 (O[13], I[13]);
  UB1DCON_14 U1 (O[14], I[14]);
endmodule

module UBCON_17_14 (O, I);
  output [17:14] O;
  input [17:14] I;
  UB1DCON_14 U0 (O[14], I[14]);
  UB1DCON_15 U1 (O[15], I[15]);
  UB1DCON_16 U2 (O[16], I[16]);
  UB1DCON_17 U3 (O[17], I[17]);
endmodule

module UBCON_19_18 (O, I);
  output [19:18] O;
  input [19:18] I;
  UB1DCON_18 U0 (O[18], I[18]);
  UB1DCON_19 U1 (O[19], I[19]);
endmodule

module UBCON_1_0 (O, I);
  output [1:0] O;
  input [1:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
endmodule

module UBCON_23_22 (O, I);
  output [23:22] O;
  input [23:22] I;
  UB1DCON_22 U0 (O[22], I[22]);
  UB1DCON_23 U1 (O[23], I[23]);
endmodule

module UBCON_24_19 (O, I);
  output [24:19] O;
  input [24:19] I;
  UB1DCON_19 U0 (O[19], I[19]);
  UB1DCON_20 U1 (O[20], I[20]);
  UB1DCON_21 U2 (O[21], I[21]);
  UB1DCON_22 U3 (O[22], I[22]);
  UB1DCON_23 U4 (O[23], I[23]);
  UB1DCON_24 U5 (O[24], I[24]);
endmodule

module UBCON_26_25 (O, I);
  output [26:25] O;
  input [26:25] I;
  UB1DCON_25 U0 (O[25], I[25]);
  UB1DCON_26 U1 (O[26], I[26]);
endmodule

module UBCON_27_25 (O, I);
  output [27:25] O;
  input [27:25] I;
  UB1DCON_25 U0 (O[25], I[25]);
  UB1DCON_26 U1 (O[26], I[26]);
  UB1DCON_27 U2 (O[27], I[27]);
endmodule

module UBCON_2_0 (O, I);
  output [2:0] O;
  input [2:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
endmodule

module UBCON_31_0 (O, I);
  output [31:0] O;
  input [31:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
  UB1DCON_9 U9 (O[9], I[9]);
  UB1DCON_10 U10 (O[10], I[10]);
  UB1DCON_11 U11 (O[11], I[11]);
  UB1DCON_12 U12 (O[12], I[12]);
  UB1DCON_13 U13 (O[13], I[13]);
  UB1DCON_14 U14 (O[14], I[14]);
  UB1DCON_15 U15 (O[15], I[15]);
  UB1DCON_16 U16 (O[16], I[16]);
  UB1DCON_17 U17 (O[17], I[17]);
  UB1DCON_18 U18 (O[18], I[18]);
  UB1DCON_19 U19 (O[19], I[19]);
  UB1DCON_20 U20 (O[20], I[20]);
  UB1DCON_21 U21 (O[21], I[21]);
  UB1DCON_22 U22 (O[22], I[22]);
  UB1DCON_23 U23 (O[23], I[23]);
  UB1DCON_24 U24 (O[24], I[24]);
  UB1DCON_25 U25 (O[25], I[25]);
  UB1DCON_26 U26 (O[26], I[26]);
  UB1DCON_27 U27 (O[27], I[27]);
  UB1DCON_28 U28 (O[28], I[28]);
  UB1DCON_29 U29 (O[29], I[29]);
  UB1DCON_30 U30 (O[30], I[30]);
  UB1DCON_31 U31 (O[31], I[31]);
endmodule

module UBCON_36_34 (O, I);
  output [36:34] O;
  input [36:34] I;
  UB1DCON_34 U0 (O[34], I[34]);
  UB1DCON_35 U1 (O[35], I[35]);
  UB1DCON_36 U2 (O[36], I[36]);
endmodule

module UBCON_39_37 (O, I);
  output [39:37] O;
  input [39:37] I;
  UB1DCON_37 U0 (O[37], I[37]);
  UB1DCON_38 U1 (O[38], I[38]);
  UB1DCON_39 U2 (O[39], I[39]);
endmodule

module UBCON_3_0 (O, I);
  output [3:0] O;
  input [3:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
endmodule

module UBCON_43_40 (O, I);
  output [43:40] O;
  input [43:40] I;
  UB1DCON_40 U0 (O[40], I[40]);
  UB1DCON_41 U1 (O[41], I[41]);
  UB1DCON_42 U2 (O[42], I[42]);
  UB1DCON_43 U3 (O[43], I[43]);
endmodule

module UBCON_49_44 (O, I);
  output [49:44] O;
  input [49:44] I;
  UB1DCON_44 U0 (O[44], I[44]);
  UB1DCON_45 U1 (O[45], I[45]);
  UB1DCON_46 U2 (O[46], I[46]);
  UB1DCON_47 U3 (O[47], I[47]);
  UB1DCON_48 U4 (O[48], I[48]);
  UB1DCON_49 U5 (O[49], I[49]);
endmodule

module UBCON_49_47 (O, I);
  output [49:47] O;
  input [49:47] I;
  UB1DCON_47 U0 (O[47], I[47]);
  UB1DCON_48 U1 (O[48], I[48]);
  UB1DCON_49 U2 (O[49], I[49]);
endmodule

module UBCON_49_48 (O, I);
  output [49:48] O;
  input [49:48] I;
  UB1DCON_48 U0 (O[48], I[48]);
  UB1DCON_49 U1 (O[49], I[49]);
endmodule

module UBCON_4_0 (O, I);
  output [4:0] O;
  input [4:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
endmodule

module UBCON_58_50 (O, I);
  output [58:50] O;
  input [58:50] I;
  UB1DCON_50 U0 (O[50], I[50]);
  UB1DCON_51 U1 (O[51], I[51]);
  UB1DCON_52 U2 (O[52], I[52]);
  UB1DCON_53 U3 (O[53], I[53]);
  UB1DCON_54 U4 (O[54], I[54]);
  UB1DCON_55 U5 (O[55], I[55]);
  UB1DCON_56 U6 (O[56], I[56]);
  UB1DCON_57 U7 (O[57], I[57]);
  UB1DCON_58 U8 (O[58], I[58]);
endmodule

module UBCON_58_54 (O, I);
  output [58:54] O;
  input [58:54] I;
  UB1DCON_54 U0 (O[54], I[54]);
  UB1DCON_55 U1 (O[55], I[55]);
  UB1DCON_56 U2 (O[56], I[56]);
  UB1DCON_57 U3 (O[57], I[57]);
  UB1DCON_58 U4 (O[58], I[58]);
endmodule

module UBCON_58_55 (O, I);
  output [58:55] O;
  input [58:55] I;
  UB1DCON_55 U0 (O[55], I[55]);
  UB1DCON_56 U1 (O[56], I[56]);
  UB1DCON_57 U2 (O[57], I[57]);
  UB1DCON_58 U3 (O[58], I[58]);
endmodule

module UBCON_58_56 (O, I);
  output [58:56] O;
  input [58:56] I;
  UB1DCON_56 U0 (O[56], I[56]);
  UB1DCON_57 U1 (O[57], I[57]);
  UB1DCON_58 U2 (O[58], I[58]);
endmodule

module UBCON_5_0 (O, I);
  output [5:0] O;
  input [5:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
endmodule

module UBCON_63_59 (O, I);
  output [63:59] O;
  input [63:59] I;
  UB1DCON_59 U0 (O[59], I[59]);
  UB1DCON_60 U1 (O[60], I[60]);
  UB1DCON_61 U2 (O[61], I[61]);
  UB1DCON_62 U3 (O[62], I[62]);
  UB1DCON_63 U4 (O[63], I[63]);
endmodule

module UBCON_63_9 (O, I);
  output [63:9] O;
  input [63:9] I;
  UB1DCON_9 U0 (O[9], I[9]);
  UB1DCON_10 U1 (O[10], I[10]);
  UB1DCON_11 U2 (O[11], I[11]);
  UB1DCON_12 U3 (O[12], I[12]);
  UB1DCON_13 U4 (O[13], I[13]);
  UB1DCON_14 U5 (O[14], I[14]);
  UB1DCON_15 U6 (O[15], I[15]);
  UB1DCON_16 U7 (O[16], I[16]);
  UB1DCON_17 U8 (O[17], I[17]);
  UB1DCON_18 U9 (O[18], I[18]);
  UB1DCON_19 U10 (O[19], I[19]);
  UB1DCON_20 U11 (O[20], I[20]);
  UB1DCON_21 U12 (O[21], I[21]);
  UB1DCON_22 U13 (O[22], I[22]);
  UB1DCON_23 U14 (O[23], I[23]);
  UB1DCON_24 U15 (O[24], I[24]);
  UB1DCON_25 U16 (O[25], I[25]);
  UB1DCON_26 U17 (O[26], I[26]);
  UB1DCON_27 U18 (O[27], I[27]);
  UB1DCON_28 U19 (O[28], I[28]);
  UB1DCON_29 U20 (O[29], I[29]);
  UB1DCON_30 U21 (O[30], I[30]);
  UB1DCON_31 U22 (O[31], I[31]);
  UB1DCON_32 U23 (O[32], I[32]);
  UB1DCON_33 U24 (O[33], I[33]);
  UB1DCON_34 U25 (O[34], I[34]);
  UB1DCON_35 U26 (O[35], I[35]);
  UB1DCON_36 U27 (O[36], I[36]);
  UB1DCON_37 U28 (O[37], I[37]);
  UB1DCON_38 U29 (O[38], I[38]);
  UB1DCON_39 U30 (O[39], I[39]);
  UB1DCON_40 U31 (O[40], I[40]);
  UB1DCON_41 U32 (O[41], I[41]);
  UB1DCON_42 U33 (O[42], I[42]);
  UB1DCON_43 U34 (O[43], I[43]);
  UB1DCON_44 U35 (O[44], I[44]);
  UB1DCON_45 U36 (O[45], I[45]);
  UB1DCON_46 U37 (O[46], I[46]);
  UB1DCON_47 U38 (O[47], I[47]);
  UB1DCON_48 U39 (O[48], I[48]);
  UB1DCON_49 U40 (O[49], I[49]);
  UB1DCON_50 U41 (O[50], I[50]);
  UB1DCON_51 U42 (O[51], I[51]);
  UB1DCON_52 U43 (O[52], I[52]);
  UB1DCON_53 U44 (O[53], I[53]);
  UB1DCON_54 U45 (O[54], I[54]);
  UB1DCON_55 U46 (O[55], I[55]);
  UB1DCON_56 U47 (O[56], I[56]);
  UB1DCON_57 U48 (O[57], I[57]);
  UB1DCON_58 U49 (O[58], I[58]);
  UB1DCON_59 U50 (O[59], I[59]);
  UB1DCON_60 U51 (O[60], I[60]);
  UB1DCON_61 U52 (O[61], I[61]);
  UB1DCON_62 U53 (O[62], I[62]);
  UB1DCON_63 U54 (O[63], I[63]);
endmodule

module UBCON_6_0 (O, I);
  output [6:0] O;
  input [6:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
endmodule

module UBCON_7_0 (O, I);
  output [7:0] O;
  input [7:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
endmodule

module UBCON_8_0 (O, I);
  output [8:0] O;
  input [8:0] I;
  UB1DCON_0 U0 (O[0], I[0]);
  UB1DCON_1 U1 (O[1], I[1]);
  UB1DCON_2 U2 (O[2], I[2]);
  UB1DCON_3 U3 (O[3], I[3]);
  UB1DCON_4 U4 (O[4], I[4]);
  UB1DCON_5 U5 (O[5], I[5]);
  UB1DCON_6 U6 (O[6], I[6]);
  UB1DCON_7 U7 (O[7], I[7]);
  UB1DCON_8 U8 (O[8], I[8]);
endmodule

module UBCON_8_7 (O, I);
  output [8:7] O;
  input [8:7] I;
  UB1DCON_7 U0 (O[7], I[7]);
  UB1DCON_8 U1 (O[8], I[8]);
endmodule

module UBExtender_63_9_6000 (O, I);
  output [64:9] O;
  input [63:9] I;
  UBCON_63_9 U0 (O[63:9], I[63:9]);
  UBZero_64_64 U1 (O[64]);
endmodule

module UBKSA_64_9_63_0 (S, X, Y);
  output [65:0] S;
  input [64:9] X;
  input [63:0] Y;
  wire [64:9] Z;
  UBExtender_63_9_6000 U0 (Z[64:9], Y[63:9]);
  UBPureKSA_64_9 U1 (S[65:9], X[64:9], Z[64:9]);
  UBCON_8_0 U2 (S[8:0], Y[8:0]);
endmodule

module UBPureKSA_64_9 (S, X, Y);
  output [65:9] S;
  input [64:9] X;
  input [64:9] Y;
  wire C;
  UBPriKSA_64_9 U0 (S, X, Y, C);
  UBZero_9_9 U1 (C);
endmodule

module UBTCCONV63_65_0 (O, I);
  output [66:0] O;
  input [65:0] I;
  UBTC1CON66_0 U0 (O[0], I[0]);
  UBTC1CON66_1 U1 (O[1], I[1]);
  UBTC1CON66_2 U2 (O[2], I[2]);
  UBTC1CON66_3 U3 (O[3], I[3]);
  UBTC1CON66_4 U4 (O[4], I[4]);
  UBTC1CON66_5 U5 (O[5], I[5]);
  UBTC1CON66_6 U6 (O[6], I[6]);
  UBTC1CON66_7 U7 (O[7], I[7]);
  UBTC1CON66_8 U8 (O[8], I[8]);
  UBTC1CON66_9 U9 (O[9], I[9]);
  UBTC1CON66_10 U10 (O[10], I[10]);
  UBTC1CON66_11 U11 (O[11], I[11]);
  UBTC1CON66_12 U12 (O[12], I[12]);
  UBTC1CON66_13 U13 (O[13], I[13]);
  UBTC1CON66_14 U14 (O[14], I[14]);
  UBTC1CON66_15 U15 (O[15], I[15]);
  UBTC1CON66_16 U16 (O[16], I[16]);
  UBTC1CON66_17 U17 (O[17], I[17]);
  UBTC1CON66_18 U18 (O[18], I[18]);
  UBTC1CON66_19 U19 (O[19], I[19]);
  UBTC1CON66_20 U20 (O[20], I[20]);
  UBTC1CON66_21 U21 (O[21], I[21]);
  UBTC1CON66_22 U22 (O[22], I[22]);
  UBTC1CON66_23 U23 (O[23], I[23]);
  UBTC1CON66_24 U24 (O[24], I[24]);
  UBTC1CON66_25 U25 (O[25], I[25]);
  UBTC1CON66_26 U26 (O[26], I[26]);
  UBTC1CON66_27 U27 (O[27], I[27]);
  UBTC1CON66_28 U28 (O[28], I[28]);
  UBTC1CON66_29 U29 (O[29], I[29]);
  UBTC1CON66_30 U30 (O[30], I[30]);
  UBTC1CON66_31 U31 (O[31], I[31]);
  UBTC1CON66_32 U32 (O[32], I[32]);
  UBTC1CON66_33 U33 (O[33], I[33]);
  UBTC1CON66_34 U34 (O[34], I[34]);
  UBTC1CON66_35 U35 (O[35], I[35]);
  UBTC1CON66_36 U36 (O[36], I[36]);
  UBTC1CON66_37 U37 (O[37], I[37]);
  UBTC1CON66_38 U38 (O[38], I[38]);
  UBTC1CON66_39 U39 (O[39], I[39]);
  UBTC1CON66_40 U40 (O[40], I[40]);
  UBTC1CON66_41 U41 (O[41], I[41]);
  UBTC1CON66_42 U42 (O[42], I[42]);
  UBTC1CON66_43 U43 (O[43], I[43]);
  UBTC1CON66_44 U44 (O[44], I[44]);
  UBTC1CON66_45 U45 (O[45], I[45]);
  UBTC1CON66_46 U46 (O[46], I[46]);
  UBTC1CON66_47 U47 (O[47], I[47]);
  UBTC1CON66_48 U48 (O[48], I[48]);
  UBTC1CON66_49 U49 (O[49], I[49]);
  UBTC1CON66_50 U50 (O[50], I[50]);
  UBTC1CON66_51 U51 (O[51], I[51]);
  UBTC1CON66_52 U52 (O[52], I[52]);
  UBTC1CON66_53 U53 (O[53], I[53]);
  UBTC1CON66_54 U54 (O[54], I[54]);
  UBTC1CON66_55 U55 (O[55], I[55]);
  UBTC1CON66_56 U56 (O[56], I[56]);
  UBTC1CON66_57 U57 (O[57], I[57]);
  UBTC1CON66_58 U58 (O[58], I[58]);
  UBTC1CON66_59 U59 (O[59], I[59]);
  UBTC1CON66_60 U60 (O[60], I[60]);
  UBTC1CON66_61 U61 (O[61], I[61]);
  UBTC1CON66_62 U62 (O[62], I[62]);
  UBTCTCONV_65_63 U63 (O[66:63], I[65:63]);
endmodule

module WLCTR_32_0_32_1_3000 (S1, S2, PP0, PP1, PP2, PP3, PP4, PP5, PP6, PP7, PP8, PP9, PP10, PP11, PP12, PP13, PP14, PP15, PP16, PP17, PP18, PP19, PP20, PP21, PP22, PP23, PP24, PP25, PP26, PP27, PP28, PP29, PP30, PP31);
  output [64:9] S1;
  output [63:0] S2;
  input [32:0] PP0;
  input [32:1] PP1;
  input [41:10] PP10;
  input [42:11] PP11;
  input [43:12] PP12;
  input [44:13] PP13;
  input [45:14] PP14;
  input [46:15] PP15;
  input [47:16] PP16;
  input [48:17] PP17;
  input [49:18] PP18;
  input [50:19] PP19;
  input [33:2] PP2;
  input [51:20] PP20;
  input [52:21] PP21;
  input [53:22] PP22;
  input [54:23] PP23;
  input [55:24] PP24;
  input [56:25] PP25;
  input [57:26] PP26;
  input [58:27] PP27;
  input [59:28] PP28;
  input [60:29] PP29;
  input [34:3] PP3;
  input [61:30] PP30;
  input [62:31] PP31;
  input [35:4] PP4;
  input [36:5] PP5;
  input [37:6] PP6;
  input [38:7] PP7;
  input [39:8] PP8;
  input [40:9] PP9;
  wire [33:2] IC0;
  wire [36:5] IC1;
  wire [55:24] IC10;
  wire [58:27] IC11;
  wire [61:30] IC12;
  wire [37:4] IC13;
  wire [44:10] IC14;
  wire [47:16] IC15;
  wire [53:20] IC16;
  wire [56:25] IC17;
  wire [62:29] IC18;
  wire [40:5] IC19;
  wire [39:8] IC2;
  wire [48:14] IC20;
  wire [54:21] IC21;
  wire [62:28] IC22;
  wire [44:6] IC23;
  wire [55:19] IC24;
  wire [63:29] IC25;
  wire [50:7] IC26;
  wire [63:26] IC27;
  wire [59:8] IC28;
  wire [42:11] IC3;
  wire [34:3] IC4;
  wire [40:7] IC5;
  wire [43:12] IC6;
  wire [46:15] IC7;
  wire [49:18] IC8;
  wire [52:21] IC9;
  wire [33:0] IS0;
  wire [36:3] IS1;
  wire [55:22] IS10;
  wire [58:25] IS11;
  wire [61:28] IS12;
  wire [39:0] IS13;
  wire [43:7] IS14;
  wire [49:13] IS15;
  wire [52:18] IS16;
  wire [58:22] IS17;
  wire [61:27] IS18;
  wire [43:0] IS19;
  wire [39:6] IS2;
  wire [49:10] IS20;
  wire [58:18] IS21;
  wire [62:25] IS22;
  wire [49:0] IS23;
  wire [58:14] IS24;
  wire [62:25] IS25;
  wire [58:0] IS26;
  wire [63:19] IS27;
  wire [63:0] IS28;
  wire [42:9] IS3;
  wire [36:0] IS4;
  wire [39:5] IS5;
  wire [43:9] IS6;
  wire [46:13] IS7;
  wire [49:16] IS8;
  wire [52:19] IS9;
  CSA_32_0_32_1_33_000 U0 (IC0, IS0, PP0, PP1, PP2);
  CSA_34_3_35_4_36_000 U1 (IC1, IS1, PP3, PP4, PP5);
  CSA_37_6_38_7_39_000 U2 (IC2, IS2, PP6, PP7, PP8);
  CSA_40_9_41_10_42000 U3 (IC3, IS3, PP9, PP10, PP11);
  CSA_33_0_33_2_36_000 U4 (IC4, IS4, IS0, IC0, IS1);
  CSA_36_5_39_6_39_000 U5 (IC5, IS5, IC1, IS2, IC2);
  CSA_42_9_42_11_43000 U6 (IC6, IS6, IS3, IC3, PP12);
  CSA_44_13_45_14_4000 U7 (IC7, IS7, PP13, PP14, PP15);
  CSA_47_16_48_17_4000 U8 (IC8, IS8, PP16, PP17, PP18);
  CSA_50_19_51_20_5000 U9 (IC9, IS9, PP19, PP20, PP21);
  CSA_53_22_54_23_5000 U10 (IC10, IS10, PP22, PP23, PP24);
  CSA_56_25_57_26_5000 U11 (IC11, IS11, PP25, PP26, PP27);
  CSA_59_28_60_29_6000 U12 (IC12, IS12, PP28, PP29, PP30);
  CSA_36_0_34_3_39_000 U13 (IC13, IS13, IS4, IC4, IS5);
  CSA_40_7_43_9_43_000 U14 (IC14, IS14, IC5, IS6, IC6);
  CSA_46_13_46_15_4000 U15 (IC15, IS15, IS7, IC7, IS8);
  CSA_49_18_52_19_5000 U16 (IC16, IS16, IC8, IS9, IC9);
  CSA_55_22_55_24_5000 U17 (IC17, IS17, IS10, IC10, IS11);
  CSA_58_27_61_28_6000 U18 (IC18, IS18, IC11, IS12, IC12);
  CSA_39_0_37_4_43_000 U19 (IC19, IS19, IS13, IC13, IS14);
  CSA_44_10_49_13_4000 U20 (IC20, IS20, IC14, IS15, IC15);
  CSA_52_18_53_20_5000 U21 (IC21, IS21, IS16, IC16, IS17);
  CSA_56_25_61_27_6000 U22 (IC22, IS22, IC17, IS18, IC18);
  CSA_43_0_40_5_49_000 U23 (IC23, IS23, IS19, IC19, IS20);
  CSA_48_14_58_18_5000 U24 (IC24, IS24, IC20, IS21, IC21);
  CSA_62_25_62_28_6000 U25 (IC25, IS25, IS22, IC22, PP31);
  CSA_49_0_44_6_58_000 U26 (IC26, IS26, IS23, IC23, IS24);
  CSA_55_19_62_25_6000 U27 (IC27, IS27, IC24, IS25, IC25);
  CSA_58_0_50_7_63_000 U28 (IC28, IS28, IS26, IC26, IS27);
  CSA_63_0_59_8_63_000 U29 (S1, S2, IS28, IC28, IC27);
endmodule

